-- MIT License
-- 
-- Copyright (c) 2019 J. Tetteroo
-- 
-- Permission is hereby granted, free of charge, to any person obtaining a copy
-- of this software and associated documentation files (the "Software"), to deal
-- in the Software without restriction, including without limitation the rights
-- to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
-- copies of the Software, and to permit persons to whom the Software is
-- furnished to do so, subject to the following conditions:
-- 
-- The above copyright notice and this permission notice shall be included in all
-- copies or substantial portions of the Software.
-- 
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
-- IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
-- FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
-- AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
-- LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
-- OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
-- SOFTWARE.

-------------------------------------------------------------------------------
--
-- Title       : tictactoe_ram
-- Design      : tictactoe
-- Author      : J. Tetteroo
-- Year		   : 2019
--
-------------------------------------------------------------------------------

-------------------------------------------------------------------------------
--
-- Description : Memory unit that stores all possible game moves in native BRAM blocks (ice40 512x8) in 3 byte records.
--
-------------------------------------------------------------------------------

library ieee;
library work;
--library ice;	-- uncomment for simulation, comment for synthesis
use ieee.std_logic_1164.all;
--use ice.vcomponent_vital.all; -- uncomment for simulation, comment for synthesis



use work.components.all; 	-- comment for simulation, uncomment for synthesis
use work.tictactoe_global.all;
use ieee.numeric_std.all;

entity tictactoe_ram is
port (
    input : in tictactoe_ram_input_type;
    output : out tictactoe_ram_output_type;
    
    clk : in std_logic;
    reset : in std_logic
    );
end tictactoe_ram;




architecture rtl of tictactoe_ram is 

	-- ### START COMMENT BLOCK FOR SYNTHESIS (comment this block when synthesizing)
	-- Component declaration of the "sb_ram512x8(sb_ram512x8_arch)" unit defined in
	-- file: "./src/sb_ice_syn_vital.vhd"
--	component sb_ram512x8
--	generic(
--		INIT_0 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
--		INIT_1 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
--		INIT_2 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
--		INIT_3 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
--		INIT_4 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
--		INIT_5 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
--		INIT_6 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
--		INIT_7 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
--		INIT_8 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
--		INIT_9 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
--		INIT_A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
--		INIT_B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
--		INIT_C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
--		INIT_D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
--		INIT_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
--		INIT_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000"
--	);
--	port(
--		RDATA : out STD_LOGIC_VECTOR(7 downto 0);
--		RCLK : in STD_LOGIC;
--		RCLKE : in STD_LOGIC := 'H';
--		RE : in STD_LOGIC := 'L';
--		RADDR : in STD_LOGIC_VECTOR(8 downto 0);
--		WCLK : in STD_LOGIC;
--		WCLKE : in STD_LOGIC := 'H';
--		WE : in STD_LOGIC := 'L';
--		WADDR : in STD_LOGIC_VECTOR(8 downto 0);
--		WDATA : in STD_LOGIC_VECTOR(7 downto 0)
--	);
--	end component;
--	for all: sb_ram512x8 use entity ice.sb_ram512x8(sb_ram512x8_arch);
	-- ### END COMMENT BLOCK FOR SYNTHESIS
    
    type t_RDATA_a is array (0 to 27) of std_logic_vector(7 downto 0);
    type t_RADDR_a is array (0 to 27) of std_logic_vector(8 downto 0);
    subtype t_RADDR is std_logic_vector(8 downto 0);
    subtype t_RCLKE is std_logic_vector(27 downto 0);
    subtype t_RE is std_logic_vector(27 downto 0);
    
    type state_type is (st_set_addr, st_wait_1, st_read_1, st_wait_2, st_read_2, st_wait_3, st_read_3, st_check, st_match, st_no_match);
    
    type reg_type is record
        match : std_logic;
        perm_block : natural range 0 to 27;      -- BRAM block
        perm_addr : natural range 0 to 511;       -- address within BRAM
		
        board_config : std_logic_vector(17 downto 0);
        output_move : std_logic_vector(3 downto 0);
        state : state_type;
	end record;
    
    signal r, rin : reg_type := (match => '0',
								perm_block => 0,
								perm_addr => 0,
								board_config => (others => '0'),
								output_move => (others => '0'),
								state => st_set_addr);
    
    signal RDATA_a : t_RDATA_a := (others => (others => '0'));
    signal RADDR_c : t_RADDR :=  (others => '0');
    signal RCLKE_c : t_RCLKE := (others => '0');
    signal RE_c : t_RE := (others => '0');
    signal RCLK_c : std_logic := '0';
    
    -- RADDR can fan out to each BRAM, we only read the relevant block, could be inefficient

begin
ram512x8_inst_0 : SB_RAM512X8
generic map (
INIT_0 => X"204000A02400802000C012008010008004002022004010004001002004000000",
INIT_1 => X"4801803001802401801301202001002401401101001001000200604000404000",
INIT_2 => X"00C08800A0800080800060800040840020840120600140540140400120400100",
INIT_3 => X"80300280200280120220200200200240110200100200000060C400A0A000C090",
INIT_4 => X"5303004303803003003303002003001302206002405102404102204002004002",
INIT_5 => X"0280920280800220A00240910240800220800200800320600300630340500300",
INIT_6 => X"A1070081000061060041000021000260C00240C00220C002A0A00280A002C092",
INIT_7 => X"1001810101212201411001410201210201010000614200A12100C11000C10800",
INIT_8 => X"04000000C18300A18300618601614201414201214201A12101812101C1100181",
INIT_9 => X"4054044041042044040042048030048020048010042024040024044012040016",
INIT_A => X"8005206005006405405405005405004405803005003405002405001404206104",
INIT_B => X"0420C004A0A00480A004C0900480900480800420A00440920440800420800400",
INIT_C => X"20600600650640500600550600450680300600350600200600150460C00440C1",
INIT_D => X"C10620C00600C10680B00680A00680920620A00600A006409206009206008006",
INIT_E => X"04C1100481100481000421210441100441000421000401000620E00640D10640",
INIT_F => X"811005212105012005411005011005010004614204414204214204A121048120"
)
port map (
RDATA => RDATA_a(0),
RADDR => RADDR_c,
RCLK => RCLK_c,
RCLKE => RCLKE_c(0),
RE => RE_c(0),
WADDR => (others => '0'),
WCLK=> '0',
WCLKE => '0',
WDATA => (others => '0'),
WE => '0'
);
ram512x8_inst_1 : SB_RAM512X8
generic map (
INIT_0 => X"8004618604418604218605216205415005414005214205014005813005812005",
INIT_1 => X"00A2000082040062060042040022020461C204A1A004C19004C18004A1800481",
INIT_2 => X"821001820201222001421001420201220201020000624000A22200C21400C200",
INIT_3 => X"0002020000C28400A28400628401624001424001224001A22201822201C21101",
INIT_4 => X"02424002224002A22002822002C2100282110282000222200242110242000222",
INIT_5 => X"2240030240038232038222038212032220030222034211030210030200026240",
INIT_6 => X"A002C29102C28002A28002828002628002428002228003226003425103424003",
INIT_7 => X"01C30801A30001830801630001430801230200C30800A3050063050262C002A2",
INIT_8 => X"803008802408801008202008002008401108001008000401634201A32201C310",
INIT_9 => X"5009004809803409003009002809001608206008405108404008204008004008",
INIT_A => X"08C0940880900880840820A00840900840840820840800800900680940500900",
INIT_B => X"40510A00570A00400A00360A00200A00160860C30840C10820C008A0A40880A0",
INIT_C => X"C00A20A00A00A00A40900A00900A00800B00680B00530B00360A20600A00680A",
INIT_D => X"0881010821210841100841030821050801000A20E00A40D10A40C10A20C00A00",
INIT_E => X"012109411009011009010808614508414008214008A12108812108C110088110",
INIT_F => X"8308818308618308418308218309415009414809014009813009812109811009"
)
port map (
RDATA => RDATA_a(1),
RADDR => RADDR_c,
RCLK => RCLK_c,
RCLKE => RCLKE_c(1),
RE => RE_c(1),
WADDR => (others => '0'),
WCLK=> '0',
WCLKE => '0',
WDATA => (others => '0'),
WE => '0'
);
ram512x8_inst_2 : SB_RAM512X8
generic map (
INIT_0 => X"0C00570C00440C80300C00360C00240C00160861C308A1A008C19008C18308A1",
INIT_1 => X"20A00C00A00C40900C00900C00800D00680D00540D00340C20600C00680C4051",
INIT_2 => X"680E00570E00360C20E00C40D10C40C00C20C00C00C00C80B00C80A00C80900C",
INIT_3 => X"0C01100C01000E20E00E00E80E40D10E00D70E00C00E00B60E00A60E00960E00",
INIT_4 => X"21610C41500C41400C21450C01400C81300C81200C81100C21210C01210C4110",
INIT_5 => X"800C21800C01800D01680D41500D01500D01480D81300D01300D01210D01100C",
INIT_6 => X"0C61C00C41C00C21C00CA1A10C81A00CC1900C81900C81800C21A10C41900C41",
INIT_7 => X"224008A22008822008C214088210088204082220084211084204082200080200",
INIT_8 => X"4009024009823009822009821409022009421009021009020808624008424008",
INIT_9 => X"0862C008A2A408C29408C28408A2840882840862840842840822840942500942",
INIT_A => X"02160A22600A42510A42400A22400A02400A22200A02200A42100A02100A0200",
INIT_B => X"A00A42900A42800A22800A02800B02680B42500B02500B02400B02360B02200B",
INIT_C => X"08C31008C30508A3050883050863050843050823050A62C00A42C00A22C00A22",
INIT_D => X"240009434009832109C31009831009830809431009430809030008634508A325",
INIT_E => X"0001240001040000644400A42000C41000C40800A40000840000640000440800",
INIT_F => X"01644001444401244401A42101842301C4100184130184000124240144140144"
)
port map (
RDATA => RDATA_a(2),
RADDR => RADDR_c,
RCLK => RCLK_c,
RCLKE => RCLKE_c(2),
RE => RE_c(2),
WADDR => (others => '0'),
WCLK=> '0',
WCLKE => '0',
WDATA => (others => '0'),
WE => '0'
);
ram512x8_inst_3 : SB_RAM512X8
generic map (
INIT_0 => X"C41102841502840002242002441102440102240002040000C48800A480006480",
INIT_1 => X"1303242003042003441003041103040302644002444002244002A42002842002",
INIT_2 => X"0264800244810224800324600344500344400324400304400384330384230384",
INIT_3 => X"650601450601250600C50000A5000065060264C002A4A002C48802A480028488",
INIT_4 => X"0004242004441004440004240004040001A52101C51001C50801A50701850001",
INIT_5 => X"05441405041005040404644004444404244404A42004842004C4100484100484",
INIT_6 => X"2480052464054454054444052444050444058430058420058410052424050420",
INIT_7 => X"200644150604150604050464C404A4A004C48804A48004848004648004448804",
INIT_8 => X"0604880624600644510644400624400604400684300684200684150624200604",
INIT_9 => X"45060425060664C00644C10624C006A4A00684A00684800624A0064481062480",
INIT_A => X"2005451005450005250005050004A52004C51004C50004A50004850004650604",
INIT_B => X"00A60000660004C58004A58004658605A52105852005C5100585100585000525",
INIT_C => X"260001664001A62001C61001C60801A60701860001660601460001260000C601",
INIT_D => X"0103260003060002664002A62002C61102C60002A60002860702660002460002",
INIT_E => X"03664003464003264003A62003862003C6110386100386000326200346110346",
INIT_F => X"202010002010401410001210000001C70801A70701670602C68102A680026680"
)
port map (
RDATA => RDATA_a(3),
RADDR => RADDR_c,
RCLK => RCLK_c,
RCLKE => RCLKE_c(3),
RE => RE_c(3),
WADDR => (others => '0'),
WCLK=> '0',
WCLKE => '0',
WDATA => (others => '0'),
WE => '0'
);
ram512x8_inst_4 : SB_RAM512X8
generic map (
INIT_0 => X"3611002011001610206010405010404410204010004010803010802010801210",
INIT_1 => X"1040921040841020841000821120601100681140541100501100401180301100",
INIT_2 => X"00201200171060C41040C01020C010A0A01080A010C0921080921080841020A0",
INIT_3 => X"9212008013006313005713003612206012006812005712004712803212003612",
INIT_4 => X"1021001001001220E01220C01200C01280B21280A21280921220A01200A01200",
INIT_5 => X"614010414010214210A12010812010C110108110108100102122104110104100",
INIT_6 => X"4011214211014211813011812011811011212211012211411011011011010010",
INIT_7 => X"10A1A310C19010C18310A1831081831061831041801021831121621141501141",
INIT_8 => X"00341420601400681440541400501400481480301400361400201400121061C0",
INIT_9 => X"C21480B01480A01480901420A01400A014409214009214008015006415005415",
INIT_A => X"1600B01600A81600921600681600571600351420E01440D21440C41420C01400",
INIT_B => X"81101421201401201441101401101401001620E01600E81600D71600C71680B2",
INIT_C => X"3015013015012615011014216214415014414014214214014214813014812014",
INIT_D => X"1421A01441901441821421801401801521621501601541501501501501401581",
INIT_E => X"42041022041002001461C21441C21421C214A1A01481A014C190148190148180",
INIT_F => X"0210624010424010224010A22210822210C21410821210820410222010421010"
)
port map (
RDATA => RDATA_a(4),
RADDR => RADDR_c,
RCLK => RCLK_c,
RCLKE => RCLKE_c(4),
RE => RE_c(4),
WADDR => (others => '0'),
WCLK=> '0',
WCLKE => '0',
WDATA => (others => '0'),
WE => '0'
);
ram512x8_inst_5 : SB_RAM512X8
generic map (
INIT_0 => X"1142401122401102401182321182221182121122221102221142141102101102",
INIT_1 => X"62C410A2A410C29410C28410A284108284106284104284102284112260114250",
INIT_2 => X"1712226012224012024012823212822212821012222012022012021012020010",
INIT_3 => X"1222A01222801202801322601302601302571302401382321302361302261302",
INIT_4 => X"C30510A3051083051063051043001023051222C012A2A01282A0128292128280",
INIT_5 => X"1011831011830211232211431011430011230211030210634010A32510C31010",
INIT_6 => X"18004018803018003018002018001011634011434011234211A32211832211C3",
INIT_7 => X"00A0184090180090180080190068190050190030182060180060184050180050",
INIT_8 => X"571A00361820E01840D01840C01820C01800C01880B01880A01880901820A018",
INIT_9 => X"1801101801001A20E01A00E01A00D01A00C01A00B01A00A01A00901A00601A00",
INIT_A => X"2160184150184140182140180140188130188120188110182120180120184110",
INIT_B => X"8018218318018019016019415019015019014019813019013019012019011018",
INIT_C => X"1861C31841C01821C018A1A31881A018C1901881901881801821A01841901841",
INIT_D => X"00E01C40D01C00D01C00C01C80B01C00B01C00A01C00901C00681C00501C0030",
INIT_E => X"501C01501C01401C81301C01301C01201C01101E00E81E00D71E00B61C20E01C",
INIT_F => X"1C21A01C01A01C41901C01901C01801D01681D01501D01301C21601C01601C41"
)
port map (
RDATA => RDATA_a(5),
RADDR => RADDR_c,
RCLK => RCLK_c,
RCLKE => RCLKE_c(5),
RE => RE_c(5),
WADDR => (others => '0'),
WCLK=> '0',
WCLKE => '0',
WDATA => (others => '0'),
WE => '0'
);
ram512x8_inst_6 : SB_RAM512X8
generic map (
INIT_0 => X"42101802101802001C21E01C41D01C41C01C21C01C01C01C81B01C81A01C8190",
INIT_1 => X"1018226018425018424018224018024018823018822018821018222018022018",
INIT_2 => X"1842841822801802801902601942501902501902401982301902301902201902",
INIT_3 => X"02101862C01842C01822C018A2A41882A018C2941882901882841822A0184290",
INIT_4 => X"901A02801B02601B02501B02361A22601A02601A02501A02401A02301A02201A",
INIT_5 => X"1823201843101843001823051803001A22E01A22C01A02C01A22A01A02A01A02",
INIT_6 => X"431019031019030018634018434018234018A32518832018C310188310188300",
INIT_7 => X"1410440410240410040419435019434019034019833019832019831019032019",
INIT_8 => X"11040310644410444410244410A42010842010C4141084151084041024201044",
INIT_9 => X"4454114444112440110444118433118420118413112420110423114414110414",
INIT_A => X"151204071064C410A4A010C48810A48010848810648010448410248311246411",
INIT_B => X"1304231304101224601224401204401284351284201284151224201204231204",
INIT_C => X"84A81284881224A0122480120487132460130463130453130440138433130433",
INIT_D => X"0610A52010C51010C50810A5071085001065061045001025061224C012A4A012",
INIT_E => X"10658611A52011852011C5101185101185001125261145101145001125061105",
INIT_F => X"044414843014842014841014242014042414441414041014040810C58810A583"
)
port map (
RDATA => RDATA_a(6),
RADDR => RADDR_c,
RCLK => RCLK_c,
RCLKE => RCLKE_c(6),
RE => RE_c(6),
WADDR => (others => '0'),
WCLK=> '0',
WCLKE => '0',
WDATA => (others => '0'),
WE => '0'
);
ram512x8_inst_7 : SB_RAM512X8
generic map (
INIT_0 => X"5415045415044415843015043415042415041414246414445414444414244414",
INIT_1 => X"1424C414A4A01484A01484881424A01444841424801404881524641504641544",
INIT_2 => X"04881624601604651604551604401684351604351604251604151464C41444C4",
INIT_3 => X"261445101445001425061405061624E01624C01604C71684A81624A01604A816",
INIT_4 => X"15252615052615451015051015050014A52014852014C5101485101485001425",
INIT_5 => X"260414A5A014C58814A580148580146586144580142586158530158520158510",
INIT_6 => X"0411260611060010664410A62010C61410C60010A60710860710660010460410",
INIT_7 => X"11664011464411264011A62011862011C6141186101186041126201146141146",
INIT_8 => X"264012A62012862012861712860712262012260012060010C68410A684106684",
INIT_9 => X"8013266013264013064013863013862013861713262013062013061713060712",
INIT_A => X"11870011670611470611270610C70810A70710670612A6A012A6801286871226",
INIT_B => X"C81000C80800A80000880000680600480000280211A72011C71011C70811A707",
INIT_C => X"2401C81001881301880401282201481001480601280201080200684000A82400",
INIT_D => X"02480002280002080000C88000A88000688001684201484001284001A8220188",
INIT_E => X"080002684002484002284002A82002882002C812028810028800022820024810",
INIT_F => X"5303484303284003084003883003882003881003282003082003481303081203"
)
port map (
RDATA => RDATA_a(7),
RADDR => RADDR_c,
RCLK => RCLK_c,
RCLKE => RCLKE_c(7),
RE => RE_c(7),
WADDR => (others => '0'),
WCLK=> '0',
WCLKE => '0',
WDATA => (others => '0'),
WE => '0'
);
ram512x8_inst_8 : SB_RAM512X8
generic map (
INIT_0 => X"0268C002A8A002C89202C88002A8800288800268800248860228800328600348",
INIT_1 => X"694201C91001C90801A90701890701690001490801290200C90000A907006902",
INIT_2 => X"4404A82004882004C81004881004880004282404481004480604280404080001",
INIT_3 => X"0588300588240588100528240508240548140508100508040468420448400428",
INIT_4 => X"C88004A880048880046886044886042880052862054854054844052840050842",
INIT_5 => X"300688200688100628200608200648150608100608000468C004A8A004C89004",
INIT_6 => X"0628A00648920648820628800608800628600648550648450628400608400688",
INIT_7 => X"69060449060429070668C00648C00628C006A8A00688A006C892068890068880",
INIT_8 => X"1005890005491005490005290205090004694204C91004C90004A90704890004",
INIT_9 => X"00CA0200AA00006A0004C98004A98004698605694205494205294205C9100589",
INIT_A => X"4A06022A00016A4001AA2201CA1001CA0801AA00018A02016A00014A08012A00",
INIT_B => X"10034A00032A00030A02026A4002AA2002CA1202CA0002AA00028A00026A0002",
INIT_C => X"026A80036A40034A40032A4003AA20038A2003CA12038A12038A02032A20034A",
INIT_D => X"880408282408481008480608280008080401CB0801AB02016B0002CA8002AA80",
INIT_E => X"2409481309081409080008684508484008284008A82408882408C81408881008",
INIT_F => X"0888800868860848860828840948500948480908430988340988240988140908"
)
port map (
RDATA => RDATA_a(8),
RADDR => RADDR_c,
RCLK => RCLK_c,
RCLKE => RCLKE_c(8),
RE => RE_c(8),
WADDR => (others => '0'),
WCLK=> '0',
WCLKE => '0',
WDATA => (others => '0'),
WE => '0'
);
ram512x8_inst_9 : SB_RAM512X8
generic map (
INIT_0 => X"08450A28200A08200A48160A08130A08000868C008A8A408C89008C88008A880",
INIT_1 => X"630B48530B08530B08400B08330B08200B08100A28600A48500A48400A28400A",
INIT_2 => X"0849080829050A68C00A48C00A28C00A28A00A48960A48860A28800A08800B08",
INIT_3 => X"891009890709491009490809090808694508C91008C90808A907088907086900",
INIT_4 => X"100C28240C08240C48140C08140C080408C98308A98708698609494809C91009",
INIT_5 => X"0D08340D08240D08140C28640C48500C48440C28450C08450C88300C88240C88",
INIT_6 => X"88800C28A40C48960C48860C28840C08860D08640D48540D08540D08400D8834",
INIT_7 => X"450E08350E08200E08100C68C00C48C00C28C00CA8A40C88A00CC8900C88900C",
INIT_8 => X"0E08C00E28A00E08A00E48960E08960E08860E28600E08650E48550E08550E08",
INIT_9 => X"C9100C89100C89000C49100C49060C29070C09070E28E00E48D00E48C00E28C0",
INIT_A => X"870D49500D49480D09480D89100D49100D09100D09070C69450C49400C29450C",
INIT_B => X"086A00084A06082A000C69C00CC9900CC9800CA9870C89800C69860C49860C29",
INIT_C => X"8A14098A00094A10094A08090A04086A4008AA2408CA1408CA0008AA00088A04",
INIT_D => X"200A4A160A4A060A2A000A0A0008CA8408AA84086A84094A48098A2409CA1409",
INIT_E => X"0B4A500B4A400B0A480B0A200B4A160B0A160B0A000A6A400A4A400A2A400A2A",
INIT_F => X"CB1009CB08098B08094B0808CB0808AB05086B050A6AC00A6A800A4A800A2A80"
)
port map (
RDATA => RDATA_a(9),
RADDR => RADDR_c,
RCLK => RCLK_c,
RCLKE => RCLKE_c(9),
RE => RE_c(9),
WADDR => (others => '0'),
WCLK=> '0',
WCLKE => '0',
WDATA => (others => '0'),
WE => '0'
);
ram512x8_inst_10 : SB_RAM512X8
generic map (
INIT_0 => X"2001CC1001CC0001AC00018C00016C00014C00012C0000CC0000AC00006C0009",
INIT_1 => X"026C4002AC2002CC1002CC0002AC00028C00026C00024C00022C00016C4001AC",
INIT_2 => X"2C4003AC20038C2003CC10038C13038C00032C20034C13034C00032C00030C00",
INIT_3 => X"00044C00042C0001CD0001AD07016D0602CC8802AC80026C80036C40034C4003",
INIT_4 => X"054C10054C00052C00050C00046C4004AC2004CC1004CC0004AC00048C00046C",
INIT_5 => X"AC80046C80056C40054C44052C4405AC20058C2005CC10058C10058C00052C24",
INIT_6 => X"20068C2006CC10068C10068C00062C20064C15064C00062C00060C0004CC8004",
INIT_7 => X"06ACA006CC8006AC80068C80066C80064C80062C80066C40064C40062C4006AC",
INIT_8 => X"CD1005CD0005AD00058D00056D00054D00052D0004CD0004AD00046D06066CC0",
INIT_9 => X"00038E00036E00034E00032E0002CE0802AE00026E0001CE0801AE00016E0005",
INIT_A => X"208011202024200022204011200012200004036E4003AE2003CE1003CE0003AE",
INIT_B => X"8031210036210024210013202061204051204041202041200041208031208021",
INIT_C => X"812020A120409220408420208420008221206121006821405121005721004821",
INIT_D => X"2200362200212200122060C42040C12020C120A0A12080A120C0922080922080",
INIT_E => X"4092220092220081230068230057230036220068224051220057220048228031",
INIT_F => X"122041032021012001012240D12240C12200C12280B22280A12280922200A122"
)
port map (
RDATA => RDATA_a(10),
RADDR => RADDR_c,
RCLK => RCLK_c,
RCLKE => RCLKE_c(10),
RE => RE_c(10),
WADDR => (others => '0'),
WCLK=> '0',
WCLKE => '0',
WDATA => (others => '0'),
WE => '0'
);
ram512x8_inst_11 : SB_RAM512X8
generic map (
INIT_0 => X"21010120614220414220214220A12120812120C1132081112081032021212041",
INIT_1 => X"4152214142212142210142218131218121218113212121210121214111210111",
INIT_2 => X"162061C120A1A320C19320C18320A18320818320618320418320218321216221",
INIT_3 => X"2500642500542500362420642400612440522400512400472400362400262400",
INIT_4 => X"00362420E12440D22440C22420C42400C22420A12400A1244092240092240086",
INIT_5 => X"112401062600E82640D22600D12600C82600B62600A126009226006826005526",
INIT_6 => X"2501212501162421612441522441422421412401422421212401212441162401",
INIT_7 => X"21A1244192244186242186240181252161250161254152250151250141250136",
INIT_8 => X"152082122082042022212042112042042022042002012461C22441C22421C224",
INIT_9 => X"21222121022221421121021121020220624420424120224120A22420822220C2",
INIT_A => X"6284204284202284212261214251214241212241210241218232218222218211",
INIT_B => X"122202212242112202112202012062C420A2A420C29120C28420A28420828420",
INIT_C => X"2302482382322302362302282302112242512242412202412282322282212282",
INIT_D => X"42C12282A122C292228292228281224291224281220281230268234251230257",
INIT_E => X"0221030220634120A32120C31520C30520A30520830520630520430520230522",
INIT_F => X"21434221234221A32121832121C3112183112183012123222143112143022123"
)
port map (
RDATA => RDATA_a(11),
RADDR => RADDR_c,
RCLK => RCLK_c,
RCLKE => RCLKE_c(11),
RE => RE_c(11),
WADDR => (others => '0'),
WCLK=> '0',
WCLKE => '0',
WDATA => (others => '0'),
WE => '0'
);
ram512x8_inst_12 : SB_RAM512X8
generic map (
INIT_0 => X"0031282061280061284051280051280041288031280031280021280011216342",
INIT_1 => X"C12880B12880A12880912820A12800A128409128009128008129006829005729",
INIT_2 => X"2A00B12A00A12A00912A00682A00572A00362820E12840D12840C12820C12800",
INIT_3 => X"81212881112821212801212841112801112801012A00E12A40D12A00D12A00C1",
INIT_4 => X"4129813129013129012129011128216128415128414128214128014128813128",
INIT_5 => X"2881912881832821A12841912841832821812801812901612941512901512901",
INIT_6 => X"00A12C00912C00612C00572C00362861C32841C12821C128A1A12881A128C193",
INIT_7 => X"212C01112E00E82E00D72E00B62C20E12C00E12C40D12C00D12C00C12C00B12C",
INIT_8 => X"2C01812D01612D01572D01312C21612C01612C41512C01512C01412C01312C01",
INIT_9 => X"02112802012C21E12C41D12C41C12C21C12C01C12C21A12C01A12C41912C0191",
INIT_A => X"6128425128424128224128024128823128822128821128222128022128421128",
INIT_B => X"2822842802812902612942512902512902412982312902312902212902112822",
INIT_C => X"62C42842C12822C128A2A42882A128C2942882912882842822A1284291284284",
INIT_D => X"812B02682B02572B02362A02612A42512A02512A02412A02312A02212A021128",
INIT_E => X"2843112843052823052803012A42D12A42C12A02C12A02A12A42912A02912A02",
INIT_F => X"031129030128634528434128234128A32128832128C315288311288301282321"
)
port map (
RDATA => RDATA_a(12),
RADDR => RADDR_c,
RCLK => RCLK_c,
RCLKE => RCLKE_c(12),
RE => RE_c(12),
WADDR => (others => '0'),
WCLK=> '0',
WCLKE => '0',
WDATA => (others => '0'),
WE => '0'
);
ram512x8_inst_13 : SB_RAM512X8
generic map (
INIT_0 => X"0820240120040329435129434129034129833129832129831129032129431129",
INIT_1 => X"20644420444420244420A42120842320C4152084132084012024232044152044",
INIT_2 => X"4444212444210444218433218423218413212424210423214413210413210403",
INIT_3 => X"082064C420A4A120C48820A48120848320648120448820248321246421445421",
INIT_4 => X"2304132244512244412204412284332284212284152204232244152204152204",
INIT_5 => X"84A3228488224488220488230463234451230453230441238433230433230421",
INIT_6 => X"0121050620A52320C51320C50120A5012085032065062045062025062244C122",
INIT_7 => X"20A58320658621A52121852321C5132185132185032125212145162145062125",
INIT_8 => X"246424445124444424244424044424242124042424441524041524040120C583",
INIT_9 => X"8624248124048625246425046425445425045425044425043425042125041124",
INIT_A => X"2644552604552604412604352604212604152464C42444C12424C42424A12444",
INIT_B => X"05062425262445162445062425062405062644C82604C82604A6260488260465",
INIT_C => X"0820660120460420260424658624458624258625252125052625451625051625",
INIT_D => X"21262421461121460421260421060120664420A62420C61520C60820A6012086",
INIT_E => X"C68820A68420668421664421464421264421A62421862121C611218611218604",
INIT_F => X"1123061123060822464122862822C61522861522860822461122460122060120"
)
port map (
RDATA => RDATA_a(13),
RADDR => RADDR_c,
RCLK => RCLK_c,
RCLKE => RCLKE_c(13),
RE => RE_c(13),
WADDR => (others => '0'),
WCLK=> '0',
WCLKE => '0',
WDATA => (others => '0'),
WE => '0'
);
ram512x8_inst_14 : SB_RAM512X8
generic map (
INIT_0 => X"22C6882286882246812346512346412306412386312386282386112306282346",
INIT_1 => X"A72121C71121C70821A70721870121670621470621270620C70820A707206706",
INIT_2 => X"5231003630206230006230405230005230004230803230003230002230001221",
INIT_3 => X"3000C23080B23080A23080923020A23000A23040923000923000823100623100",
INIT_4 => X"80B23200B23200A23200923200683200573200323020E23040D23040C23020C2",
INIT_5 => X"323081223081123021223001223041123001123001023200E23200D23200C232",
INIT_6 => X"3101423181323101323101223101123021623041523041423021423001423081",
INIT_7 => X"81923081833021A2304192304182302182300182312162310162314152310152",
INIT_8 => X"A23400923400623400523400363061C23041C23021C230A1A33081A230C19230",
INIT_9 => X"3401123600E83600D23600B23420E23400E23440D23400D23400C23400B23400",
INIT_A => X"0182350162350152350136342162340162344152340152340142340132340122",
INIT_B => X"123002023421E23441D23441C23421C23401C23421A23401A234419234019234",
INIT_C => X"3042523042423022423002423082323082223082123022223002223042123002",
INIT_D => X"0282312262310262314252310252310242318232310232310222310212302262",
INIT_E => X"C23022C230A2A43082A230C2923082923082823022A230429230428430228430",
INIT_F => X"3302573302363202623202523202423282323202323202223202123062C43042"
)
port map (
RDATA => RDATA_a(14),
RADDR => RADDR_c,
RCLK => RCLK_c,
RCLKE => RCLKE_c(14),
RE => RE_c(14),
WADDR => (others => '0'),
WCLK=> '0',
WCLKE => '0',
WDATA => (others => '0'),
WE => '0'
);
ram512x8_inst_15 : SB_RAM512X8
generic map (
INIT_0 => X"43023023023003023202C23282B23282A23282923202A2320292320282330268",
INIT_1 => X"0230634230434230234230A32530832230C31530831230830530232230431230",
INIT_2 => X"3143423123423103423183323183223183123123223103223143123103123103",
INIT_3 => X"0444308433308423308415302424300426304414300413300405312362314352",
INIT_4 => X"5431045331044431843331043631042631041630246430445430444430244430",
INIT_5 => X"3024C430A4A33084A33084833024A33044843024843004833124643104633144",
INIT_6 => X"04573304363204683204573204433284353204333204283204153064C43044C4",
INIT_7 => X"033025263045133045033025033005063204C73284A83204A832048833046833",
INIT_8 => X"31851331252631052631451631051631050630A52330852330C5153085133085",
INIT_9 => X"042634041530A5A330C58330A583308583306583304583302583318533318523",
INIT_A => X"A634048635046435045435043634246434046434445434045434044434043634",
INIT_B => X"3604C83604A83604683604553604353424E43444C43424C43404C43424A43404",
INIT_C => X"25863405863505363505263505163425263405263445153405163405063604E8",
INIT_D => X"2430C6153086153086053026243046143046043026043006043425A634458634",
INIT_E => X"31861431262431062431461431061431060430664430464430264430A6243086",
INIT_F => X"8684306684304684302684312664314654314644312644310644318634318624"
)
port map (
RDATA => RDATA_a(15),
RADDR => RADDR_c,
RCLK => RCLK_c,
RCLKE => RCLKE_c(15),
RE => RE_c(15),
WADDR => (others => '0'),
WCLK=> '0',
WCLKE => '0',
WDATA => (others => '0'),
WE => '0'
);
ram512x8_inst_16 : SB_RAM512X8
generic map (
INIT_0 => X"453286353286283286153206283206173206053066C430A6A430C68430A68430",
INIT_1 => X"3027053286A83286883206873306683306573306473306363306283306173206",
INIT_2 => X"471631470631270631070630A72530C71530C70530A705308705306705304705",
INIT_3 => X"1220880220282420481220480620280420080331872831871731870731272631",
INIT_4 => X"21082421481321081321080420684420484220284220A82420882320C8132088",
INIT_5 => X"4886202883212862214852214844212842210844218833218824218813212824",
INIT_6 => X"222248122208132208022068C420A8A320C89220C88220A88220888220688220",
INIT_7 => X"2388322308332308222308132248522248482208432288322288222288122208",
INIT_8 => X"88A222C892228892228882224892224888220882230863234853230853230842",
INIT_9 => X"0221090720694220C91320C90220A9072089032069062049062029072248C822",
INIT_A => X"20A98320698621694221494221294221C9132189132189072149122149062129",
INIT_B => X"286424485224484424284424084424282424082424481624081424080220C983",
INIT_C => X"8624288224088425286425086425485425085425084425083425082425081224",
INIT_D => X"2608552608422608352608222608122468C42448C22428C42428A42448962448",
INIT_E => X"29062409062648D22648C82608C82608A2264892260896260882260865264855",
INIT_F => X"4225294225094225491625091625090624694224494224294224491624490624"
)
port map (
RDATA => RDATA_a(16),
RADDR => RADDR_c,
RCLK => RCLK_c,
RCLKE => RCLKE_c(16),
RE => RE_c(16),
WADDR => (others => '0'),
WCLK=> '0',
WCLKE => '0',
WDATA => (others => '0'),
WE => '0'
);
ram512x8_inst_17 : SB_RAM512X8
generic map (
INIT_0 => X"20AA02208A04206A02204A08202A022469C22469862449862429862549522549",
INIT_1 => X"8A12218A04212A22214A12214A08212A02210A08206A4220AA2420CA1220CA08",
INIT_2 => X"08220A0220CA8420AA84206A84216A42214A48212A4221AA24218A2421CA1221",
INIT_3 => X"230A22234A12230A12230A08224A48228A2222CA12228A12228A02224A12224A",
INIT_4 => X"6B0522CA9222CA82228A82224A82234A52234A48230A48238A32238A22238A12",
INIT_5 => X"04216B4221CB1221CB0821AB07218B07216B02214B08212B0220CB0820AB0720",
INIT_6 => X"2848442828432808482888332888242888132828242808242848132808162808",
INIT_7 => X"0884290868294853290857290848298834290833290824290817282864284853",
INIT_8 => X"C32828C428A8A42888A328C8932888932888832828A428489628488428288428",
INIT_9 => X"2B08572B08362A08682A48532A08572A08482A08362A08232A08162868C42848",
INIT_A => X"49032829052809072A48D32A48C82A08C82A08A32A48962A08962A08832B0868",
INIT_B => X"1729491329091729090728694528494328294528C91328891328890328491328",
INIT_C => X"28C99328C98328A9832889832869832849832829832949532949482909482989",
INIT_D => X"08572D08342C28642C08642C48542C08572C08472C08362C08242C08162869C3",
INIT_E => X"E42C48D42C48C42C28C42C08C42C28A42C08A42C48962C08962C08862D08642D",
INIT_F => X"2C09072E08E82E08D72E08C82E08B62E08A62E08962E08682E08572E08362C28"
)
port map (
RDATA => RDATA_a(17),
RADDR => RADDR_c,
RCLK => RCLK_c,
RCLKE => RCLKE_c(17),
RE => RE_c(17),
WADDR => (others => '0'),
WCLK=> '0',
WCLKE => '0',
WDATA => (others => '0'),
WE => '0'
);
ram512x8_inst_18 : SB_RAM512X8
generic map (
INIT_0 => X"29872C09862D09572D09472D09172C49552C49452C29472C09472C49162C0916",
INIT_1 => X"14288A04282A24284A14284A04282A04280A042C49C82C29C72C49962C49862C",
INIT_2 => X"290A24294A14290A14290A08286A44284A48282A4428AA24288A2428CA14288A",
INIT_3 => X"AA84288A84286A84284A84282A84294A54294A48290A48298A34298A24298A14",
INIT_4 => X"552A4A482A0A482A0A252A4A162A0A162A0A05286AC428AAA428CA9428CA8428",
INIT_5 => X"2A4AC82A4A962A4A862A0A862B0A682B0A572B0A482B0A362B0A262B0A162A4A",
INIT_6 => X"4B16294B08290B08286B4528CB1528CB0528AB05288B05286B05284B05282B05",
INIT_7 => X"2320CC1320CC0320AC03208C03206C03204C03202C03294B48298B17298B0729",
INIT_8 => X"218C2321CC13218C13218C03212C24214C13214C03212C04210C03206C4420AC",
INIT_9 => X"8C03224C15224C08220C0320CC8320AC83206C83216C44214C44212C4421AC24",
INIT_A => X"33238C23238C13230C23234C13230C13230C03224C43228C2322CC15228C1322",
INIT_B => X"212D0320CD0320AD03206D0622CC88228C83224C88234C53234C43230C43238C",
INIT_C => X"2C24244C15244C04242C04240C0421CD1321CD0321AD07218D03216D06214D06",
INIT_D => X"44252C44250C44252C24250C24254C14250C14250C04246C44244C44242C4424",
INIT_E => X"260C25264C15260C15260C05246CC4246C84244C86242C84252C64254C54254C",
INIT_F => X"2D06250D06246D06244D06242D06264CC8264C88260C86264C55264C45260C45"
)
port map (
RDATA => RDATA_a(18),
RADDR => RADDR_c,
RCLK => RCLK_c,
RCLKE => RCLKE_c(18),
RE => RE_c(18),
WADDR => (others => '0'),
WCLK=> '0',
WCLKE => '0',
WDATA => (others => '0'),
WE => '0'
);
ram512x8_inst_19 : SB_RAM512X8
generic map (
INIT_0 => X"04218E08216E04214E08212E0420CE0820AE04206E04246D86254D16254D0625",
INIT_1 => X"234E08230E0822CE1522CE08228E08224E08216E4421AE2421CE1421CE0821AE",
INIT_2 => X"500600300221CF0821AF07216F0622CE88234E48238E28238E17238E08234E16",
INIT_3 => X"1401500201300201100200704100B02200D01400D00100B00100900200700600",
INIT_4 => X"00708101704201504101304201B02201902201D0110190140190020130220150",
INIT_5 => X"902202D01102901102900202302202501102500102300202100100D08100B082",
INIT_6 => X"2103901103302103102203501103101103100302704102504102304302B02202",
INIT_7 => X"0290810270810250810230860330620350510350430330430310430390310390",
INIT_8 => X"710101510801310200D10800B1020071020270C102B0A202D09102D08102B081",
INIT_9 => X"0104302504501404500204300204100101714201B12201D10801B10101910801",
INIT_A => X"05501405101405100404704204504404304504B02104902404D0110490140490",
INIT_B => X"3081053061055054055044053041051042059034059024059014053021051022",
INIT_C => X"110610110610050470C104B0A104D09104D08804B08704908204708604508104",
INIT_D => X"0630650650510650410630450610410690310690210690110630250610220650",
INIT_E => X"30C106B0A20690A206D0920690920690820630A1065091065081063081061081",
INIT_F => X"0104714204B12104D10804B1070491080471060451080431010670C10650C106"
)
port map (
RDATA => RDATA_a(19),
RADDR => RADDR_c,
RCLK => RCLK_c,
RCLKE => RCLKE_c(19),
RE => RE_c(19),
WADDR => (others => '0'),
WCLK=> '0',
WCLKE => '0',
WDATA => (others => '0'),
WE => '0'
);
ram512x8_inst_20 : SB_RAM512X8
generic map (
INIT_0 => X"04718605714205514105314205B1210591210591010531220551010531020511",
INIT_1 => X"D20101B20101920101720601520601320200D20100B20100720604D18804B187",
INIT_2 => X"0602B22202D21102D20102B20102920102720602520102320601B22201D21401",
INIT_3 => X"02728103B22203922203D2110392110392020332220352110352010332020312",
INIT_4 => X"900108302408501408500608300108100501D30801B30101730202D28102B281",
INIT_5 => X"2309501309101409100108704308504308304508B02108902408D01408901408",
INIT_6 => X"0890840870860850840830860950510950430910430990340990210990140910",
INIT_7 => X"10430A30210A10230A50110A10110A10060870C308B0A408D09408D08108B081",
INIT_8 => X"630B50530B10530B10430B10330B10210B10110A30650A50510A50430A30430A",
INIT_9 => X"0851080831050A70C30A50C10A30C30A30A60A50910A50810A30860A10810B10",
INIT_A => X"514809912809910809510809110808714508B12508D10808B101089108087101",
INIT_B => X"340C90240C90140C30250C10240C50140C10140C100408D18808B18708718609",
INIT_C => X"0D10410D90340D10340D10210D10140C30650C50540C50440C30450C10450C90",
INIT_D => X"D0940C90940C90840C30A10C50940C50840C30840C10810D10640D50540D1054",
INIT_E => X"510E10550E10450E10350E10210E10110C70C10C50C10C30C10CB0A40C90A40C",
INIT_F => X"0E50C10E30C10E10C10E30A60E10A60E50910E10910E10860E30650E10650E50"
)
port map (
RDATA => RDATA_a(20),
RADDR => RADDR_c,
RCLK => RCLK_c,
RCLKE => RCLKE_c(20),
RE => RE_c(20),
WADDR => (others => '0'),
WCLK=> '0',
WCLKE => '0',
WDATA => (others => '0'),
WE => '0'
);
ram512x8_inst_21 : SB_RAM512X8
generic map (
INIT_0 => X"51480C31450CB1210C91210C91010C31250C51080C31050C11080E30E10E50D1",
INIT_1 => X"870C91880C71860C51880C31810D51480D11480D91210D11280D11080C71450C",
INIT_2 => X"08D21408D20108B2010892040872060852060832050C71C10CB1A10CD1880CB1",
INIT_3 => X"D28408B28408728609922109D21409921409920109521109520609120608B221",
INIT_4 => X"810A32860B12260B52160B12160B12060A32250A52110A52060A32060A120608",
INIT_5 => X"00D40100B40700740109D30809930809530808D30808B3050873050A72860A52",
INIT_6 => X"540102340101744101B42101D41101D40101B401019401017401015401013401",
INIT_7 => X"1103540103340103140102744102B42102D41102D40102B40102940102740102",
INIT_8 => X"02748103744103544103344303B42103942303D4110394110394010334230354",
INIT_9 => X"D40104B40104940104740104540104340101D50801B50701750602D48102B487",
INIT_A => X"1105941405940105342405541405540105340105140404744104B42104D41104",
INIT_B => X"06340106140104D48804B48704748105744105544405344405B42105942405D4",
INIT_C => X"744106544106344106B42106942506D411069415069401063425065411065401",
INIT_D => X"0804B5070475060674C106B4A106D48106B48106948106748106548106348106",
INIT_E => X"01D60101B60701760605B52105D50105B50105950105750105550105350104D5",
INIT_F => X"B62103D61103D60103B60103960103760103560103360102D60102B607027601"
)
port map (
RDATA => RDATA_a(21),
RADDR => RADDR_c,
RCLK => RCLK_c,
RCLKE => RCLKE_c(21),
RE => RE_c(21),
WADDR => (others => '0'),
WCLK=> '0',
WCLKE => '0',
WDATA => (others => '0'),
WE => '0'
);
ram512x8_inst_22 : SB_RAM512X8
generic map (
INIT_0 => X"4310B02210902210D01410901410900410302210501410500410300410100303",
INIT_1 => X"1190341190221190141130221110231150141110141110061070431050441030",
INIT_2 => X"D08210B087109084107082105084103087113062115054115043113042111042",
INIT_3 => X"431290321290221290121230221210231210121210071070C410B0A210D09410",
INIT_4 => X"1330631310631310531310431390321310331310231310121230631230431210",
INIT_5 => X"71061051021031021230C712B0A21290A21290921290821230A2123087121082",
INIT_6 => X"2811910811312211510211310211110810714210B12210D10810B10710910810",
INIT_7 => X"14501414101414100410D18810B18710718611714211514211314211B1221191",
INIT_8 => X"1014143065145054145044143044141044149034149022149012143022141024",
INIT_9 => X"8414308414108215306215106415505415105415104415903415103415102415",
INIT_A => X"1470C41450C41430C214B0A21490A214D0921490921490881430A21450941450",
INIT_B => X"10A2161092161087163065161065161055161042169032161035161025161012",
INIT_C => X"221451021431021411081630E21630C71610C71690B21690A21690921630A216",
INIT_D => X"15912815312215112815110214714214514214314214B1221491281491081431",
INIT_E => X"B1A214D18814B187149188147186145188143182153162155142153142151142",
INIT_F => X"0611120610B22210D21410D20210B2021092041072061052041032061471C214"
)
port map (
RDATA => RDATA_a(22),
RADDR => RADDR_c,
RCLK => RCLK_c,
RCLKE => RCLKE_c(22),
RE => RE_c(22),
WADDR => (others => '0'),
WCLK=> '0',
WCLKE => '0',
WDATA => (others => '0'),
WE => '0'
);
ram512x8_inst_23 : SB_RAM512X8
generic map (
INIT_0 => X"10B28410728411B22211922211D2141192141192021132221152141152041132",
INIT_1 => X"122613121613120612B22212922212921212920212322612320612120610D284",
INIT_2 => X"0810B30510730612B2A212B28212928212328613923213922213921213322613",
INIT_3 => X"18501418101418100311B32211D30811B30211930811730611530211330210D3",
INIT_4 => X"1013183065185054185043183043181043189034189024189014183025181026",
INIT_5 => X"9418508418308318108419106819505319105319104319903419103319102819",
INIT_6 => X"1A10131870C31850C41830C318B0A41890A418D0941890941890841830A31850",
INIT_7 => X"10931A10831B10631B10531B10361A30631A10631A10571A10431A10361A1026",
INIT_8 => X"281891031831251851031831051811081A30E31A30C31A10C71A30A61A10A61A",
INIT_9 => X"18318319514319114819912819112819110818714318514318314518B1251891",
INIT_A => X"90341C10341C10281C10141871C318B1A318D18318B183189183187183185183",
INIT_B => X"941C10941C10841D10681D10541D10341C30651C10681C50541C10541C10481C",
INIT_C => X"1C30E41C50D41C50C41C30C41C10C41C90B41C90A41C90941C30A41C10A41C50",
INIT_D => X"11281C11081E10E81E10D71E10C71E10B61E10A61E10961E10681E10571E1036",
INIT_E => X"861C11881D11681D11481D11281C31651C51481C31451C11481C91281C31251C",
INIT_F => X"1852141852041832051812041C51C81C31C71C91A81C91881C31A61C51881C31"
)
port map (
RDATA => RDATA_a(23),
RADDR => RADDR_c,
RCLK => RCLK_c,
RCLKE => RCLKE_c(23),
RE => RE_c(23),
WADDR => (others => '0'),
WCLK=> '0',
WCLKE => '0',
WDATA => (others => '0'),
WE => '0'
);
ram512x8_inst_24 : SB_RAM512X8
generic map (
INIT_0 => X"921419122619521419121419120618B22418922418D214189214189204183225",
INIT_1 => X"0618B2A418D29418D28418B28418928418728418528418328419923419922419",
INIT_2 => X"1833051A32A61A32861A12861B12361B12261B12161A32261A12261A12161A12",
INIT_3 => X"340719932819930819530619130818B32518D30518B305189305187305185305",
INIT_4 => X"0411340611140410744410B42310D41410D40310B40710940710740310540410",
INIT_5 => X"11744311544411344311B42311942311D4141194141194041134231154141154",
INIT_6 => X"344312B42312942312941512940712342312340712140310D48410B487107483",
INIT_7 => X"8713346313344313144313943313942313941313342313142313141313140312",
INIT_8 => X"11950811750611550311350610D50810B50710750612B4A312B4871294871234",
INIT_9 => X"D41414941414940814342414541414540414340414140411B52311D50811B507",
INIT_A => X"1415342415142415541415141415140414744414544414344414B42414942414",
INIT_B => X"1474841454841434871534641554541554441534441514441594341594241594",
INIT_C => X"94251694151634251614251614151614051474C414B4A414D48814B487149488",
INIT_D => X"061634C71694A81694881634A616348716148716346516344516144516943516",
INIT_E => X"15352615550615350615150614B52514D50814B5071495081475061455051435",
INIT_F => X"760611560411360610D60410B60710760414D58814B587147586159528159508"
)
port map (
RDATA => RDATA_a(24),
RADDR => RADDR_c,
RCLK => RCLK_c,
RCLKE => RCLKE_c(24),
RE => RE_c(24),
WADDR => (others => '0'),
WCLK=> '0',
WCLKE => '0',
WDATA => (others => '0'),
WE => '0'
);
ram512x8_inst_25 : SB_RAM512X8
generic map (
INIT_0 => X"0613160712B62512B60712960712360711B62411D61411D60411B60711960711",
INIT_1 => X"00B80200780211D70811B70711770612B6871396281396171396071336261336",
INIT_2 => X"380201784201B82201D81201D80201B80201980201780201580201380200D802",
INIT_3 => X"0203380203180202784202B82202D81202D80202B80202980202780202580202",
INIT_4 => X"03784203584303384203B82203982203D8120398120398020338220358120358",
INIT_5 => X"B80204980204780204580204380201D90801B90201790202D88202B882027886",
INIT_6 => X"1405980205382205581405580205380205180204784204B82204D81204D80204",
INIT_7 => X"06180204D88204B88204788605784205584205384205B82205982405D8120598",
INIT_8 => X"584506384506B82206982206D812069812069802063822065812065802063802",
INIT_9 => X"020678C206B8A206D89206D88206B88206988206788206588206388206784206",
INIT_A => X"017A0205794205D90205B90205990205790205590205390204D90804B9070479",
INIT_B => X"DA0203BA02039A02037A02035A02033A0202DA0202BA02027A0601DA0201BA02",
INIT_C => X"4508B82408D81408D80308B80308980408780308580308380303BA2203DA1203",
INIT_D => X"08B88308788609584309982409D8140998140998030958140958030918030878",
INIT_E => X"18130B18030A78430A58430A38450A38230A58130A58060A38030A180308D883",
INIT_F => X"050879030A78C30A78860A58860A38860B58530B58430B18430B18230B58130B"
)
port map (
RDATA => RDATA_a(25),
RADDR => RADDR_c,
RCLK => RCLK_c,
RCLKE => RCLKE_c(25),
RE => RE_c(25),
WADDR => (others => '0'),
WCLK=> '0',
WCLKE => '0',
WDATA => (others => '0'),
WE => '0'
);
ram512x8_inst_26 : SB_RAM512X8
generic map (
INIT_0 => X"0C98040C38240C58140C58040C38040C180409D90809990809590808D90808B9",
INIT_1 => X"18240D58140D18140D18040C78450C58450C38450CB8240C98240CD8140C9814",
INIT_2 => X"840C98840C78860C58860C38860D58540D58440D18440D98340D98240D98140D",
INIT_3 => X"0E18450E38250E18250E58150E18150E18050C78C40CB8A40CD8940CD8840CB8",
INIT_4 => X"58C80E38C70E38A60E58960E58860E38860E18860E38650E58550E58450E3845",
INIT_5 => X"480D99070D59080D19080C79450CD9080CB9070C99050C79050C59080C39050E",
INIT_6 => X"09DA1409DA04099A04095A0608DA0408BA04087A050CD9880CB9870C79860D59",
INIT_7 => X"000000000000000009DB080A7A860B5A160B5A060B1A060A7A060A5A060A3A05",
INIT_8 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_9 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_F => X"0000000000000000000000000000000000000000000000000000000000000000"
)
port map (
RDATA => RDATA_a(26),
RADDR => RADDR_c,
RCLK => RCLK_c,
RCLKE => RCLKE_c(26),
RE => RE_c(26),
WADDR => (others => '0'),
WCLK=> '0',
WCLKE => '0',
WDATA => (others => '0'),
WE => '0'
);
    combinatorial : process(reset, r, RDATA_a)
	    variable v : reg_type;
    
        variable block_addr : natural range 0 to 14508; -- NUM_RECORDS=4836*3
        variable block_select : natural range 0 to 27;  -- NUM_BLOCKS
        variable block_idx : natural range 0 to 511;    -- BLOCK_SIZE
        variable block_buf : std_logic_vector(7 downto 0);
    
        begin
            v := r;
            
            block_addr := input.perm_idx * 3;
            block_select := block_addr / 512;   -- synthesizer bitshift
            block_idx := block_addr mod 512;
        
            case (r.state) is
                when st_set_addr =>
					v.board_config := "000000000000000000";
                    v.perm_block := block_select;
                    v.perm_addr := block_idx;
					
                    v.state := st_read_1;
                when st_read_1 =>
					v.board_config := "00000000000000" & RDATA_a(r.perm_block)(7 downto 4);
					--v.board_config := "0000000000" & RDATA_a(r.perm_block);
					v.output_move := RDATA_a(r.perm_block)(3 downto 0);
					
					v.perm_addr := (r.perm_addr + 1) mod 512;
				    if r.perm_addr = 511 then
                        v.perm_block := r.perm_block + 1;
                  	end if;
					  
                    v.state := st_read_2;
                when st_read_2 =>
					v.board_config := "000000" & RDATA_a(r.perm_block) & r.board_config(3 downto 0);
					--v.board_config := "0000000000" & RDATA_a(r.perm_block);
					
					v.perm_addr := (r.perm_addr + 1) mod 512;
				    if r.perm_addr = 511 then
                        v.perm_block := r.perm_block + 1;
                  	end if;
                    v.state := st_read_3;
                when st_read_3 =>
					v.board_config := RDATA_a(r.perm_block)(5 downto 0) & r.board_config(11 downto 0);
					--v.board_config := "0000000000" & RDATA_a(r.perm_block);
					
                    
                    v.state := st_check;
                when st_check =>					
                    if (v.board_config = (input.board_p1 & input.board_p2)) then
                        v.state := st_match;
                    else
                        v.state := st_no_match;
                    end if;
					
                when st_match =>
					v.state := st_match;
				
                when st_no_match =>
					v.state := st_no_match;
				when others =>
					v.state := st_set_addr;
                
                    
            end case;
			
			if (reset = '1') then
				v.state := st_set_addr;
			end if;
            
            RADDR_c <= std_logic_vector(to_unsigned(v.perm_addr, 9));
			
            RCLKE_c <= (others => '0');
            RCLKE_c(v.perm_block) <= '1';
			RCLKE_c(v.perm_block+1) <= '1';	-- enable the next block in case it overlaps, easiest but not optimal solution
			
            RE_c <= (others => '0');
            RE_c(v.perm_block) <= '1';
			RE_c(v.perm_block+1) <= '1';
			
            
            output.match <= '1' when (r.state = st_match) else '0';
            output.done <= '1' when (r.state = st_match OR r.state = st_no_match) else '0';
            output.output_move <= r.output_move;
			rin <= v;
            
    end process;

	synchronous : process(clk)
	begin
		if clk'event and clk = '1' then
			r <= rin;
		end if;
	end process;  
	
	RCLK_c <= clk;
    
end rtl;