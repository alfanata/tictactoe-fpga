-- MIT License
-- 
-- Copyright (c) 2019 J. Tetteroo
-- 
-- Permission is hereby granted, free of charge, to any person obtaining a copy
-- of this software and associated documentation files (the "Software"), to deal
-- in the Software without restriction, including without limitation the rights
-- to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
-- copies of the Software, and to permit persons to whom the Software is
-- furnished to do so, subject to the following conditions:
-- 
-- The above copyright notice and this permission notice shall be included in all
-- copies or substantial portions of the Software.
-- 
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
-- IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
-- FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
-- AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
-- LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
-- OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
-- SOFTWARE.

-------------------------------------------------------------------------------
--
-- Title       : tictactoe_ram_tb
-- Design      : tictactoe
-- Author      : J. Tetteroo
-- Year		   : 2019
--
-------------------------------------------------------------------------------

-------------------------------------------------------------------------------
--
-- Description : testbench for tictactoe_ram entity, tests all valid board configurations
--
-------------------------------------------------------------------------------

library ieee;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.tictactoe_global.all;
use work.tictactoe_ram;


entity tictactoe_ram_tb is
end tictactoe_ram_tb;


architecture test of tictactoe_ram_tb is

    constant DELTA : time := 100 ns;


    signal sim_finished : boolean := false;

    signal clk : std_logic;
    signal reset : std_logic;

    
    signal ram_input : tictactoe_ram_input_type;

    signal ram_output : tictactoe_ram_output_type;


begin
    -- ram instance
    tttram : entity tictactoe_ram
        port map(clk => clk,
                reset => reset,
                input => ram_input,
                output => ram_output);
          
    -- Test
    clock : process
    begin
        if not sim_finished then
            clk <= '1';
            wait for DELTA / 2;
            clk <= '0';
            wait for DELTA / 2;
        else
            wait;
        end if;
    end process clock;
    
    
    simulation : process
	
		procedure check_mem(constant rec_in: in natural;
							constant board_p1 : in std_logic_vector(8 downto 0);
							constant board_p2 : in std_logic_vector(8 downto 0);
							constant next_move : in natural;
							constant is_match : in std_logic) is
			variable output_move : natural;
		begin
			-- state set_addr
			ram_input.perm_idx <= rec_in;
			ram_input.board_p1 <= board_p1;
			ram_input.board_p2 <= board_p2;
			
			wait until rising_edge(clk);
			-- state read 1
			assert ram_output.done = '0' report "Operation completed prematurely" severity error;
			
        	wait until rising_edge(clk);
			-- state read 2
			assert ram_output.done = '0' report "Operation completed prematurely" severity error;
			
			wait until rising_edge(clk);
			-- state read 3
			assert ram_output.done = '0' report "Operation completed prematurely" severity error;
			
			
			wait until rising_edge(clk);
			-- state check
			assert ram_output.done = '0' report "Operation completed prematurely" severity error;
			
			-- state match/no_match
        	wait until rising_edge(clk);
			wait for DELTA / 4;
			output_move := to_integer(unsigned(ram_output.output_move));
			assert ram_output.done = '1' report "Operation not completed: " & integer'image(rec_in) severity error;
			assert ram_output.match = is_match report "Match signal mismatch: " & integer'image(rec_in) severity error;
			assert output_move = next_move report "Incorrect output move: " & integer'image(rec_in) severity error;
			
		end procedure;
		
		procedure sync_reset is
		begin
			wait until rising_edge(CLK);
			wait for DELTA / 4;
			reset <= '1';
			wait until rising_edge(CLK);
			wait for DELTA / 4;
			reset <= '0';
		end procedure sync_reset;

		variable init_input : tictactoe_ram_input_type;
    begin
		
		init_input.perm_idx := 0;
		init_input.board_p1 := "000000000";
		init_input.board_p2 := "000000000";

		ram_input <= init_input;
		reset <= '0';
		
        wait for DELTA;
		
		report "#### START TESTS ####";
sync_reset;
check_mem(0,"000000000","000000000",0,'1'); -- (0, 0, 0, 0, 0, 0, 0, 0, 0)
sync_reset;
check_mem(1,"000000001","000000000",4,'1'); -- (0, 0, 0, 0, 0, 0, 0, 0, 1)
sync_reset;
check_mem(2,"000000010","000000000",1,'1'); -- (0, 0, 0, 0, 0, 0, 0, 1, 0)
sync_reset;
check_mem(3,"000000010","000000001",0,'1'); -- (0, 0, 0, 0, 0, 0, 0, 1, 2)
sync_reset;
check_mem(4,"000000001","000000010",2,'1'); -- (0, 0, 0, 0, 0, 0, 0, 2, 1)
sync_reset;
check_mem(5,"000000100","000000000",4,'1'); -- (0, 0, 0, 0, 0, 0, 1, 0, 0)
sync_reset;
check_mem(6,"000000100","000000001",0,'1'); -- (0, 0, 0, 0, 0, 0, 1, 0, 2)
sync_reset;
check_mem(7,"000000110","000000001",2,'1'); -- (0, 0, 0, 0, 0, 0, 1, 1, 2)
sync_reset;
check_mem(8,"000000100","000000010",0,'1'); -- (0, 0, 0, 0, 0, 0, 1, 2, 0)
sync_reset;
check_mem(9,"000000101","000000010",4,'1'); -- (0, 0, 0, 0, 0, 0, 1, 2, 1)
sync_reset;
check_mem(10,"000000001","000000100",0,'1'); -- (0, 0, 0, 0, 0, 0, 2, 0, 1)
sync_reset;
check_mem(11,"000000010","000000100",0,'1'); -- (0, 0, 0, 0, 0, 0, 2, 1, 0)
sync_reset;
check_mem(12,"000000011","000000100",0,'1'); -- (0, 0, 0, 0, 0, 0, 2, 1, 1)
sync_reset;
check_mem(13,"000001000","000000000",2,'1'); -- (0, 0, 0, 0, 0, 1, 0, 0, 0)
sync_reset;
check_mem(14,"000001000","000000001",0,'1'); -- (0, 0, 0, 0, 0, 1, 0, 0, 2)
sync_reset;
check_mem(15,"000001010","000000001",1,'1'); -- (0, 0, 0, 0, 0, 1, 0, 1, 2)
sync_reset;
check_mem(16,"000001000","000000010",4,'1'); -- (0, 0, 0, 0, 0, 1, 0, 2, 0)
sync_reset;
check_mem(17,"000001001","000000010",0,'1'); -- (0, 0, 0, 0, 0, 1, 0, 2, 1)
sync_reset;
check_mem(18,"000001100","000000001",3,'1'); -- (0, 0, 0, 0, 0, 1, 1, 0, 2)
sync_reset;
check_mem(19,"000001100","000000010",4,'1'); -- (0, 0, 0, 0, 0, 1, 1, 2, 0)
sync_reset;
check_mem(20,"000001100","000000011",0,'1'); -- (0, 0, 0, 0, 0, 1, 1, 2, 2)
sync_reset;
check_mem(21,"000001000","000000100",8,'1'); -- (0, 0, 0, 0, 0, 1, 2, 0, 0)
sync_reset;
check_mem(22,"000001001","000000100",0,'1'); -- (0, 0, 0, 0, 0, 1, 2, 0, 1)
sync_reset;
check_mem(23,"000001010","000000100",0,'1'); -- (0, 0, 0, 0, 0, 1, 2, 1, 0)
sync_reset;
check_mem(24,"000001010","000000101",4,'1'); -- (0, 0, 0, 0, 0, 1, 2, 1, 2)
sync_reset;
check_mem(25,"000001001","000000110",0,'1'); -- (0, 0, 0, 0, 0, 1, 2, 2, 1)
sync_reset;
check_mem(26,"000000001","000001000",4,'1'); -- (0, 0, 0, 0, 0, 2, 0, 0, 1)
sync_reset;
check_mem(27,"000000010","000001000",4,'1'); -- (0, 0, 0, 0, 0, 2, 0, 1, 0)
sync_reset;
check_mem(28,"000000011","000001000",0,'1'); -- (0, 0, 0, 0, 0, 2, 0, 1, 1)
sync_reset;
check_mem(29,"000000100","000001000",0,'1'); -- (0, 0, 0, 0, 0, 2, 1, 0, 0)
sync_reset;
check_mem(30,"000000101","000001000",0,'1'); -- (0, 0, 0, 0, 0, 2, 1, 0, 1)
sync_reset;
check_mem(31,"000000110","000001000",8,'1'); -- (0, 0, 0, 0, 0, 2, 1, 1, 0)
sync_reset;
check_mem(32,"000000110","000001001",0,'1'); -- (0, 0, 0, 0, 0, 2, 1, 1, 2)
sync_reset;
check_mem(33,"000000101","000001010",0,'1'); -- (0, 0, 0, 0, 0, 2, 1, 2, 1)
sync_reset;
check_mem(34,"000000011","000001100",4,'1'); -- (0, 0, 0, 0, 0, 2, 2, 1, 1)
sync_reset;
check_mem(35,"000010000","000000000",0,'1'); -- (0, 0, 0, 0, 1, 0, 0, 0, 0)
sync_reset;
check_mem(36,"000010000","000000001",0,'1'); -- (0, 0, 0, 0, 1, 0, 0, 0, 2)
sync_reset;
check_mem(37,"000010010","000000001",1,'1'); -- (0, 0, 0, 0, 1, 0, 0, 1, 2)
sync_reset;
check_mem(38,"000010000","000000010",0,'1'); -- (0, 0, 0, 0, 1, 0, 0, 2, 0)
sync_reset;
check_mem(39,"000010001","000000010",0,'1'); -- (0, 0, 0, 0, 1, 0, 0, 2, 1)
sync_reset;
check_mem(40,"000010100","000000001",2,'1'); -- (0, 0, 0, 0, 1, 0, 1, 0, 2)
sync_reset;
check_mem(41,"000010100","000000010",0,'1'); -- (0, 0, 0, 0, 1, 0, 1, 2, 0)
sync_reset;
check_mem(42,"000010100","000000011",0,'1'); -- (0, 0, 0, 0, 1, 0, 1, 2, 2)
sync_reset;
check_mem(43,"000010000","000000100",0,'1'); -- (0, 0, 0, 0, 1, 0, 2, 0, 0)
sync_reset;
check_mem(44,"000010001","000000100",0,'1'); -- (0, 0, 0, 0, 1, 0, 2, 0, 1)
sync_reset;
check_mem(45,"000010010","000000100",1,'1'); -- (0, 0, 0, 0, 1, 0, 2, 1, 0)
sync_reset;
check_mem(46,"000010010","000000101",1,'1'); -- (0, 0, 0, 0, 1, 0, 2, 1, 2)
sync_reset;
check_mem(47,"000010001","000000110",0,'1'); -- (0, 0, 0, 0, 1, 0, 2, 2, 1)
sync_reset;
check_mem(48,"000011000","000000001",3,'1'); -- (0, 0, 0, 0, 1, 1, 0, 0, 2)
sync_reset;
check_mem(49,"000011000","000000010",0,'1'); -- (0, 0, 0, 0, 1, 1, 0, 2, 0)
sync_reset;
check_mem(50,"000011000","000000011",3,'1'); -- (0, 0, 0, 0, 1, 1, 0, 2, 2)
sync_reset;
check_mem(51,"000011100","000000011",0,'1'); -- (0, 0, 0, 0, 1, 1, 1, 2, 2)
sync_reset;
check_mem(52,"000011000","000000100",3,'1'); -- (0, 0, 0, 0, 1, 1, 2, 0, 0)
sync_reset;
check_mem(53,"000011000","000000101",3,'1'); -- (0, 0, 0, 0, 1, 1, 2, 0, 2)
sync_reset;
check_mem(54,"000011010","000000101",0,'1'); -- (0, 0, 0, 0, 1, 1, 2, 1, 2)
sync_reset;
check_mem(55,"000011000","000000110",3,'1'); -- (0, 0, 0, 0, 1, 1, 2, 2, 0)
sync_reset;
check_mem(56,"000011001","000000110",0,'1'); -- (0, 0, 0, 0, 1, 1, 2, 2, 1)
sync_reset;
check_mem(57,"000010000","000001000",0,'1'); -- (0, 0, 0, 0, 1, 2, 0, 0, 0)
sync_reset;
check_mem(58,"000010001","000001000",0,'1'); -- (0, 0, 0, 0, 1, 2, 0, 0, 1)
sync_reset;
check_mem(59,"000010010","000001000",0,'1'); -- (0, 0, 0, 0, 1, 2, 0, 1, 0)
sync_reset;
check_mem(60,"000010010","000001001",1,'1'); -- (0, 0, 0, 0, 1, 2, 0, 1, 2)
sync_reset;
check_mem(61,"000010001","000001010",0,'1'); -- (0, 0, 0, 0, 1, 2, 0, 2, 1)
sync_reset;
check_mem(62,"000010100","000001000",0,'1'); -- (0, 0, 0, 0, 1, 2, 1, 0, 0)
sync_reset;
check_mem(63,"000010100","000001001",2,'1'); -- (0, 0, 0, 0, 1, 2, 1, 0, 2)
sync_reset;
check_mem(64,"000010110","000001001",2,'1'); -- (0, 0, 0, 0, 1, 2, 1, 1, 2)
sync_reset;
check_mem(65,"000010100","000001010",0,'1'); -- (0, 0, 0, 0, 1, 2, 1, 2, 0)
sync_reset;
check_mem(66,"000010101","000001010",0,'1'); -- (0, 0, 0, 0, 1, 2, 1, 2, 1)
sync_reset;
check_mem(67,"000010001","000001100",0,'1'); -- (0, 0, 0, 0, 1, 2, 2, 0, 1)
sync_reset;
check_mem(68,"000010010","000001100",0,'1'); -- (0, 0, 0, 0, 1, 2, 2, 1, 0)
sync_reset;
check_mem(69,"000010011","000001100",0,'1'); -- (0, 0, 0, 0, 1, 2, 2, 1, 1)
sync_reset;
check_mem(70,"000000001","000010000",0,'1'); -- (0, 0, 0, 0, 2, 0, 0, 0, 1)
sync_reset;
check_mem(71,"000000010","000010000",0,'1'); -- (0, 0, 0, 0, 2, 0, 0, 1, 0)
sync_reset;
check_mem(72,"000000011","000010000",6,'1'); -- (0, 0, 0, 0, 2, 0, 0, 1, 1)
sync_reset;
check_mem(73,"000000100","000010000",0,'1'); -- (0, 0, 0, 0, 2, 0, 1, 0, 0)
sync_reset;
check_mem(74,"000000101","000010000",7,'1'); -- (0, 0, 0, 0, 2, 0, 1, 0, 1)
sync_reset;
check_mem(75,"000000110","000010000",8,'1'); -- (0, 0, 0, 0, 2, 0, 1, 1, 0)
sync_reset;
check_mem(76,"000000110","000010001",0,'1'); -- (0, 0, 0, 0, 2, 0, 1, 1, 2)
sync_reset;
check_mem(77,"000000101","000010010",1,'1'); -- (0, 0, 0, 0, 2, 0, 1, 2, 1)
sync_reset;
check_mem(78,"000000011","000010100",2,'1'); -- (0, 0, 0, 0, 2, 0, 2, 1, 1)
sync_reset;
check_mem(79,"000001000","000010000",0,'1'); -- (0, 0, 0, 0, 2, 1, 0, 0, 0)
sync_reset;
check_mem(80,"000001001","000010000",2,'1'); -- (0, 0, 0, 0, 2, 1, 0, 0, 1)
sync_reset;
check_mem(81,"000001010","000010000",2,'1'); -- (0, 0, 0, 0, 2, 1, 0, 1, 0)
sync_reset;
check_mem(82,"000001010","000010001",0,'1'); -- (0, 0, 0, 0, 2, 1, 0, 1, 2)
sync_reset;
check_mem(83,"000001001","000010010",2,'1'); -- (0, 0, 0, 0, 2, 1, 0, 2, 1)
sync_reset;
check_mem(84,"000001100","000010000",1,'1'); -- (0, 0, 0, 0, 2, 1, 1, 0, 0)
sync_reset;
check_mem(85,"000001100","000010001",0,'1'); -- (0, 0, 0, 0, 2, 1, 1, 0, 2)
sync_reset;
check_mem(86,"000001110","000010001",0,'1'); -- (0, 0, 0, 0, 2, 1, 1, 1, 2)
sync_reset;
check_mem(87,"000001100","000010010",1,'1'); -- (0, 0, 0, 0, 2, 1, 1, 2, 0)
sync_reset;
check_mem(88,"000001101","000010010",1,'1'); -- (0, 0, 0, 0, 2, 1, 1, 2, 1)
sync_reset;
check_mem(89,"000001001","000010100",2,'1'); -- (0, 0, 0, 0, 2, 1, 2, 0, 1)
sync_reset;
check_mem(90,"000001010","000010100",2,'1'); -- (0, 0, 0, 0, 2, 1, 2, 1, 0)
sync_reset;
check_mem(91,"000001011","000010100",2,'1'); -- (0, 0, 0, 0, 2, 1, 2, 1, 1)
sync_reset;
check_mem(92,"000000011","000011000",6,'1'); -- (0, 0, 0, 0, 2, 2, 0, 1, 1)
sync_reset;
check_mem(93,"000000101","000011000",3,'1'); -- (0, 0, 0, 0, 2, 2, 1, 0, 1)
sync_reset;
check_mem(94,"000000110","000011000",3,'1'); -- (0, 0, 0, 0, 2, 2, 1, 1, 0)
sync_reset;
check_mem(95,"000100000","000000000",0,'1'); -- (0, 0, 0, 1, 0, 0, 0, 0, 0)
sync_reset;
check_mem(96,"000100000","000000001",6,'1'); -- (0, 0, 0, 1, 0, 0, 0, 0, 2)
sync_reset;
check_mem(97,"000100010","000000001",2,'1'); -- (0, 0, 0, 1, 0, 0, 0, 1, 2)
sync_reset;
check_mem(98,"000100000","000000010",4,'1'); -- (0, 0, 0, 1, 0, 0, 0, 2, 0)
sync_reset;
check_mem(99,"000100001","000000010",4,'1'); -- (0, 0, 0, 1, 0, 0, 0, 2, 1)
sync_reset;
check_mem(100,"000100100","000000001",0,'1'); -- (0, 0, 0, 1, 0, 0, 1, 0, 2)
sync_reset;
check_mem(101,"000100100","000000010",0,'1'); -- (0, 0, 0, 1, 0, 0, 1, 2, 0)
sync_reset;
check_mem(102,"000100100","000000011",0,'1'); -- (0, 0, 0, 1, 0, 0, 1, 2, 2)
sync_reset;
check_mem(103,"000100000","000000100",2,'1'); -- (0, 0, 0, 1, 0, 0, 2, 0, 0)
sync_reset;
check_mem(104,"000100001","000000100",4,'1'); -- (0, 0, 0, 1, 0, 0, 2, 0, 1)
sync_reset;
check_mem(105,"000100010","000000100",1,'1'); -- (0, 0, 0, 1, 0, 0, 2, 1, 0)
sync_reset;
check_mem(106,"000100010","000000101",4,'1'); -- (0, 0, 0, 1, 0, 0, 2, 1, 2)
sync_reset;
check_mem(107,"000100001","000000110",1,'1'); -- (0, 0, 0, 1, 0, 0, 2, 2, 1)
sync_reset;
check_mem(108,"000101000","000000001",4,'1'); -- (0, 0, 0, 1, 0, 1, 0, 0, 2)
sync_reset;
check_mem(109,"000101000","000000010",4,'1'); -- (0, 0, 0, 1, 0, 1, 0, 2, 0)
sync_reset;
check_mem(110,"000101000","000000011",4,'1'); -- (0, 0, 0, 1, 0, 1, 0, 2, 2)
sync_reset;
check_mem(111,"000101100","000000011",0,'1'); -- (0, 0, 0, 1, 0, 1, 1, 2, 2)
sync_reset;
check_mem(112,"000101000","000000100",4,'1'); -- (0, 0, 0, 1, 0, 1, 2, 0, 0)
sync_reset;
check_mem(113,"000101000","000000101",4,'1'); -- (0, 0, 0, 1, 0, 1, 2, 0, 2)
sync_reset;
check_mem(114,"000101010","000000101",4,'1'); -- (0, 0, 0, 1, 0, 1, 2, 1, 2)
sync_reset;
check_mem(115,"000101000","000000110",4,'1'); -- (0, 0, 0, 1, 0, 1, 2, 2, 0)
sync_reset;
check_mem(116,"000101001","000000110",0,'1'); -- (0, 0, 0, 1, 0, 1, 2, 2, 1)
sync_reset;
check_mem(117,"000100000","000001000",0,'1'); -- (0, 0, 0, 1, 0, 2, 0, 0, 0)
sync_reset;
check_mem(118,"000100001","000001000",0,'1'); -- (0, 0, 0, 1, 0, 2, 0, 0, 1)
sync_reset;
check_mem(119,"000100010","000001000",0,'1'); -- (0, 0, 0, 1, 0, 2, 0, 1, 0)
sync_reset;
check_mem(120,"000100010","000001001",2,'1'); -- (0, 0, 0, 1, 0, 2, 0, 1, 2)
sync_reset;
check_mem(121,"000100001","000001010",0,'1'); -- (0, 0, 0, 1, 0, 2, 0, 2, 1)
sync_reset;
check_mem(122,"000100100","000001000",0,'1'); -- (0, 0, 0, 1, 0, 2, 1, 0, 0)
sync_reset;
check_mem(123,"000100100","000001001",0,'1'); -- (0, 0, 0, 1, 0, 2, 1, 0, 2)
sync_reset;
check_mem(124,"000100110","000001001",0,'1'); -- (0, 0, 0, 1, 0, 2, 1, 1, 2)
sync_reset;
check_mem(125,"000100100","000001010",0,'1'); -- (0, 0, 0, 1, 0, 2, 1, 2, 0)
sync_reset;
check_mem(126,"000100101","000001010",0,'1'); -- (0, 0, 0, 1, 0, 2, 1, 2, 1)
sync_reset;
check_mem(127,"000100001","000001100",0,'1'); -- (0, 0, 0, 1, 0, 2, 2, 0, 1)
sync_reset;
check_mem(128,"000100010","000001100",1,'1'); -- (0, 0, 0, 1, 0, 2, 2, 1, 0)
sync_reset;
check_mem(129,"000100011","000001100",0,'1'); -- (0, 0, 0, 1, 0, 2, 2, 1, 1)
sync_reset;
check_mem(130,"000110000","000000001",5,'1'); -- (0, 0, 0, 1, 1, 0, 0, 0, 2)
sync_reset;
check_mem(131,"000110000","000000010",0,'1'); -- (0, 0, 0, 1, 1, 0, 0, 2, 0)
sync_reset;
check_mem(132,"000110000","000000011",5,'1'); -- (0, 0, 0, 1, 1, 0, 0, 2, 2)
sync_reset;
check_mem(133,"000110100","000000011",0,'1'); -- (0, 0, 0, 1, 1, 0, 1, 2, 2)
sync_reset;
check_mem(134,"000110000","000000100",5,'1'); -- (0, 0, 0, 1, 1, 0, 2, 0, 0)
sync_reset;
check_mem(135,"000110000","000000101",5,'1'); -- (0, 0, 0, 1, 1, 0, 2, 0, 2)
sync_reset;
check_mem(136,"000110010","000000101",0,'1'); -- (0, 0, 0, 1, 1, 0, 2, 1, 2)
sync_reset;
check_mem(137,"000110000","000000110",5,'1'); -- (0, 0, 0, 1, 1, 0, 2, 2, 0)
sync_reset;
check_mem(138,"000110001","000000110",0,'1'); -- (0, 0, 0, 1, 1, 0, 2, 2, 1)
sync_reset;
check_mem(139,"000110000","000001000",0,'1'); -- (0, 0, 0, 1, 1, 2, 0, 0, 0)
sync_reset;
check_mem(140,"000110000","000001001",2,'1'); -- (0, 0, 0, 1, 1, 2, 0, 0, 2)
sync_reset;
check_mem(141,"000110010","000001001",2,'1'); -- (0, 0, 0, 1, 1, 2, 0, 1, 2)
sync_reset;
check_mem(142,"000110000","000001010",0,'1'); -- (0, 0, 0, 1, 1, 2, 0, 2, 0)
sync_reset;
check_mem(143,"000110001","000001010",0,'1'); -- (0, 0, 0, 1, 1, 2, 0, 2, 1)
sync_reset;
check_mem(144,"000110100","000001001",2,'1'); -- (0, 0, 0, 1, 1, 2, 1, 0, 2)
sync_reset;
check_mem(145,"000110100","000001010",0,'1'); -- (0, 0, 0, 1, 1, 2, 1, 2, 0)
sync_reset;
check_mem(146,"000110100","000001011",0,'1'); -- (0, 0, 0, 1, 1, 2, 1, 2, 2)
sync_reset;
check_mem(147,"000110000","000001100",1,'1'); -- (0, 0, 0, 1, 1, 2, 2, 0, 0)
sync_reset;
check_mem(148,"000110001","000001100",0,'1'); -- (0, 0, 0, 1, 1, 2, 2, 0, 1)
sync_reset;
check_mem(149,"000110010","000001100",1,'1'); -- (0, 0, 0, 1, 1, 2, 2, 1, 0)
sync_reset;
check_mem(150,"000110010","000001101",1,'1'); -- (0, 0, 0, 1, 1, 2, 2, 1, 2)
sync_reset;
check_mem(151,"000110001","000001110",0,'1'); -- (0, 0, 0, 1, 1, 2, 2, 2, 1)
sync_reset;
check_mem(152,"000100000","000010000",0,'1'); -- (0, 0, 0, 1, 2, 0, 0, 0, 0)
sync_reset;
check_mem(153,"000100001","000010000",0,'1'); -- (0, 0, 0, 1, 2, 0, 0, 0, 1)
sync_reset;
check_mem(154,"000100010","000010000",0,'1'); -- (0, 0, 0, 1, 2, 0, 0, 1, 0)
sync_reset;
check_mem(155,"000100010","000010001",0,'1'); -- (0, 0, 0, 1, 2, 0, 0, 1, 2)
sync_reset;
check_mem(156,"000100001","000010010",1,'1'); -- (0, 0, 0, 1, 2, 0, 0, 2, 1)
sync_reset;
check_mem(157,"000100100","000010000",0,'1'); -- (0, 0, 0, 1, 2, 0, 1, 0, 0)
sync_reset;
check_mem(158,"000100100","000010001",0,'1'); -- (0, 0, 0, 1, 2, 0, 1, 0, 2)
sync_reset;
check_mem(159,"000100110","000010001",0,'1'); -- (0, 0, 0, 1, 2, 0, 1, 1, 2)
sync_reset;
check_mem(160,"000100100","000010010",0,'1'); -- (0, 0, 0, 1, 2, 0, 1, 2, 0)
sync_reset;
check_mem(161,"000100101","000010010",1,'1'); -- (0, 0, 0, 1, 2, 0, 1, 2, 1)
sync_reset;
check_mem(162,"000100001","000010100",2,'1'); -- (0, 0, 0, 1, 2, 0, 2, 0, 1)
sync_reset;
check_mem(163,"000100010","000010100",2,'1'); -- (0, 0, 0, 1, 2, 0, 2, 1, 0)
sync_reset;
check_mem(164,"000100011","000010100",2,'1'); -- (0, 0, 0, 1, 2, 0, 2, 1, 1)
sync_reset;
check_mem(165,"000101000","000010000",0,'1'); -- (0, 0, 0, 1, 2, 1, 0, 0, 0)
sync_reset;
check_mem(166,"000101000","000010001",0,'1'); -- (0, 0, 0, 1, 2, 1, 0, 0, 2)
sync_reset;
check_mem(167,"000101010","000010001",0,'1'); -- (0, 0, 0, 1, 2, 1, 0, 1, 2)
sync_reset;
check_mem(168,"000101000","000010010",0,'1'); -- (0, 0, 0, 1, 2, 1, 0, 2, 0)
sync_reset;
check_mem(169,"000101001","000010010",1,'1'); -- (0, 0, 0, 1, 2, 1, 0, 2, 1)
sync_reset;
check_mem(170,"000101100","000010001",0,'1'); -- (0, 0, 0, 1, 2, 1, 1, 0, 2)
sync_reset;
check_mem(171,"000101100","000010010",0,'1'); -- (0, 0, 0, 1, 2, 1, 1, 2, 0)
sync_reset;
check_mem(172,"000101100","000010011",0,'1'); -- (0, 0, 0, 1, 2, 1, 1, 2, 2)
sync_reset;
check_mem(173,"000101000","000010100",0,'1'); -- (0, 0, 0, 1, 2, 1, 2, 0, 0)
sync_reset;
check_mem(174,"000101001","000010100",2,'1'); -- (0, 0, 0, 1, 2, 1, 2, 0, 1)
sync_reset;
check_mem(175,"000101010","000010100",0,'1'); -- (0, 0, 0, 1, 2, 1, 2, 1, 0)
sync_reset;
check_mem(176,"000101010","000010101",0,'1'); -- (0, 0, 0, 1, 2, 1, 2, 1, 2)
sync_reset;
check_mem(177,"000101001","000010110",2,'1'); -- (0, 0, 0, 1, 2, 1, 2, 2, 1)
sync_reset;
check_mem(178,"000100001","000011000",6,'1'); -- (0, 0, 0, 1, 2, 2, 0, 0, 1)
sync_reset;
check_mem(179,"000100010","000011000",6,'1'); -- (0, 0, 0, 1, 2, 2, 0, 1, 0)
sync_reset;
check_mem(180,"000100011","000011000",6,'1'); -- (0, 0, 0, 1, 2, 2, 0, 1, 1)
sync_reset;
check_mem(181,"000100100","000011000",0,'1'); -- (0, 0, 0, 1, 2, 2, 1, 0, 0)
sync_reset;
check_mem(182,"000100101","000011000",0,'1'); -- (0, 0, 0, 1, 2, 2, 1, 0, 1)
sync_reset;
check_mem(183,"000100110","000011000",0,'1'); -- (0, 0, 0, 1, 2, 2, 1, 1, 0)
sync_reset;
check_mem(184,"000100110","000011001",0,'1'); -- (0, 0, 0, 1, 2, 2, 1, 1, 2)
sync_reset;
check_mem(185,"000100101","000011010",0,'1'); -- (0, 0, 0, 1, 2, 2, 1, 2, 1)
sync_reset;
check_mem(186,"000100011","000011100",2,'1'); -- (0, 0, 0, 1, 2, 2, 2, 1, 1)
sync_reset;
check_mem(187,"000000001","000100000",2,'1'); -- (0, 0, 0, 2, 0, 0, 0, 0, 1)
sync_reset;
check_mem(188,"000000010","000100000",4,'1'); -- (0, 0, 0, 2, 0, 0, 0, 1, 0)
sync_reset;
check_mem(189,"000000011","000100000",6,'1'); -- (0, 0, 0, 2, 0, 0, 0, 1, 1)
sync_reset;
check_mem(190,"000000100","000100000",4,'1'); -- (0, 0, 0, 2, 0, 0, 1, 0, 0)
sync_reset;
check_mem(191,"000000101","000100000",0,'1'); -- (0, 0, 0, 2, 0, 0, 1, 0, 1)
sync_reset;
check_mem(192,"000000110","000100000",0,'1'); -- (0, 0, 0, 2, 0, 0, 1, 1, 0)
sync_reset;
check_mem(193,"000000110","000100001",4,'1'); -- (0, 0, 0, 2, 0, 0, 1, 1, 2)
sync_reset;
check_mem(194,"000000101","000100010",2,'1'); -- (0, 0, 0, 2, 0, 0, 1, 2, 1)
sync_reset;
check_mem(195,"000000011","000100100",0,'1'); -- (0, 0, 0, 2, 0, 0, 2, 1, 1)
sync_reset;
check_mem(196,"000001000","000100000",0,'1'); -- (0, 0, 0, 2, 0, 1, 0, 0, 0)
sync_reset;
check_mem(197,"000001001","000100000",2,'1'); -- (0, 0, 0, 2, 0, 1, 0, 0, 1)
sync_reset;
check_mem(198,"000001010","000100000",2,'1'); -- (0, 0, 0, 2, 0, 1, 0, 1, 0)
sync_reset;
check_mem(199,"000001010","000100001",0,'1'); -- (0, 0, 0, 2, 0, 1, 0, 1, 2)
sync_reset;
check_mem(200,"000001001","000100010",0,'1'); -- (0, 0, 0, 2, 0, 1, 0, 2, 1)
sync_reset;
check_mem(201,"000001100","000100000",2,'1'); -- (0, 0, 0, 2, 0, 1, 1, 0, 0)
sync_reset;
check_mem(202,"000001100","000100001",0,'1'); -- (0, 0, 0, 2, 0, 1, 1, 0, 2)
sync_reset;
check_mem(203,"000001110","000100001",1,'1'); -- (0, 0, 0, 2, 0, 1, 1, 1, 2)
sync_reset;
check_mem(204,"000001100","000100010",2,'1'); -- (0, 0, 0, 2, 0, 1, 1, 2, 0)
sync_reset;
check_mem(205,"000001101","000100010",2,'1'); -- (0, 0, 0, 2, 0, 1, 1, 2, 1)
sync_reset;
check_mem(206,"000001001","000100100",0,'1'); -- (0, 0, 0, 2, 0, 1, 2, 0, 1)
sync_reset;
check_mem(207,"000001010","000100100",0,'1'); -- (0, 0, 0, 2, 0, 1, 2, 1, 0)
sync_reset;
check_mem(208,"000001011","000100100",0,'1'); -- (0, 0, 0, 2, 0, 1, 2, 1, 1)
sync_reset;
check_mem(209,"000000011","000101000",4,'1'); -- (0, 0, 0, 2, 0, 2, 0, 1, 1)
sync_reset;
check_mem(210,"000000101","000101000",4,'1'); -- (0, 0, 0, 2, 0, 2, 1, 0, 1)
sync_reset;
check_mem(211,"000000110","000101000",4,'1'); -- (0, 0, 0, 2, 0, 2, 1, 1, 0)
sync_reset;
check_mem(212,"000010000","000100000",0,'1'); -- (0, 0, 0, 2, 1, 0, 0, 0, 0)
sync_reset;
check_mem(213,"000010001","000100000",0,'1'); -- (0, 0, 0, 2, 1, 0, 0, 0, 1)
sync_reset;
check_mem(214,"000010010","000100000",0,'1'); -- (0, 0, 0, 2, 1, 0, 0, 1, 0)
sync_reset;
check_mem(215,"000010010","000100001",1,'1'); -- (0, 0, 0, 2, 1, 0, 0, 1, 2)
sync_reset;
check_mem(216,"000010001","000100010",0,'1'); -- (0, 0, 0, 2, 1, 0, 0, 2, 1)
sync_reset;
check_mem(217,"000010100","000100000",0,'1'); -- (0, 0, 0, 2, 1, 0, 1, 0, 0)
sync_reset;
check_mem(218,"000010100","000100001",1,'1'); -- (0, 0, 0, 2, 1, 0, 1, 0, 2)
sync_reset;
check_mem(219,"000010110","000100001",0,'1'); -- (0, 0, 0, 2, 1, 0, 1, 1, 2)
sync_reset;
check_mem(220,"000010100","000100010",0,'1'); -- (0, 0, 0, 2, 1, 0, 1, 2, 0)
sync_reset;
check_mem(221,"000010101","000100010",0,'1'); -- (0, 0, 0, 2, 1, 0, 1, 2, 1)
sync_reset;
check_mem(222,"000010001","000100100",0,'1'); -- (0, 0, 0, 2, 1, 0, 2, 0, 1)
sync_reset;
check_mem(223,"000010010","000100100",0,'1'); -- (0, 0, 0, 2, 1, 0, 2, 1, 0)
sync_reset;
check_mem(224,"000010011","000100100",0,'1'); -- (0, 0, 0, 2, 1, 0, 2, 1, 1)
sync_reset;
check_mem(225,"000011000","000100000",0,'1'); -- (0, 0, 0, 2, 1, 1, 0, 0, 0)
sync_reset;
check_mem(226,"000011000","000100001",0,'1'); -- (0, 0, 0, 2, 1, 1, 0, 0, 2)
sync_reset;
check_mem(227,"000011010","000100001",1,'1'); -- (0, 0, 0, 2, 1, 1, 0, 1, 2)
sync_reset;
check_mem(228,"000011000","000100010",2,'1'); -- (0, 0, 0, 2, 1, 1, 0, 2, 0)
sync_reset;
check_mem(229,"000011001","000100010",0,'1'); -- (0, 0, 0, 2, 1, 1, 0, 2, 1)
sync_reset;
check_mem(230,"000011100","000100001",2,'1'); -- (0, 0, 0, 2, 1, 1, 1, 0, 2)
sync_reset;
check_mem(231,"000011100","000100010",2,'1'); -- (0, 0, 0, 2, 1, 1, 1, 2, 0)
sync_reset;
check_mem(232,"000011100","000100011",2,'1'); -- (0, 0, 0, 2, 1, 1, 1, 2, 2)
sync_reset;
check_mem(233,"000011000","000100100",0,'1'); -- (0, 0, 0, 2, 1, 1, 2, 0, 0)
sync_reset;
check_mem(234,"000011001","000100100",0,'1'); -- (0, 0, 0, 2, 1, 1, 2, 0, 1)
sync_reset;
check_mem(235,"000011010","000100100",0,'1'); -- (0, 0, 0, 2, 1, 1, 2, 1, 0)
sync_reset;
check_mem(236,"000011010","000100101",1,'1'); -- (0, 0, 0, 2, 1, 1, 2, 1, 2)
sync_reset;
check_mem(237,"000011001","000100110",0,'1'); -- (0, 0, 0, 2, 1, 1, 2, 2, 1)
sync_reset;
check_mem(238,"000010001","000101000",0,'1'); -- (0, 0, 0, 2, 1, 2, 0, 0, 1)
sync_reset;
check_mem(239,"000010010","000101000",0,'1'); -- (0, 0, 0, 2, 1, 2, 0, 1, 0)
sync_reset;
check_mem(240,"000010011","000101000",0,'1'); -- (0, 0, 0, 2, 1, 2, 0, 1, 1)
sync_reset;
check_mem(241,"000010100","000101000",0,'1'); -- (0, 0, 0, 2, 1, 2, 1, 0, 0)
sync_reset;
check_mem(242,"000010101","000101000",0,'1'); -- (0, 0, 0, 2, 1, 2, 1, 0, 1)
sync_reset;
check_mem(243,"000010110","000101000",0,'1'); -- (0, 0, 0, 2, 1, 2, 1, 1, 0)
sync_reset;
check_mem(244,"000010110","000101001",1,'1'); -- (0, 0, 0, 2, 1, 2, 1, 1, 2)
sync_reset;
check_mem(245,"000010101","000101010",0,'1'); -- (0, 0, 0, 2, 1, 2, 1, 2, 1)
sync_reset;
check_mem(246,"000010011","000101100",0,'1'); -- (0, 0, 0, 2, 1, 2, 2, 1, 1)
sync_reset;
check_mem(247,"000000011","000110000",5,'1'); -- (0, 0, 0, 2, 2, 0, 0, 1, 1)
sync_reset;
check_mem(248,"000000101","000110000",5,'1'); -- (0, 0, 0, 2, 2, 0, 1, 0, 1)
sync_reset;
check_mem(249,"000000110","000110000",8,'1'); -- (0, 0, 0, 2, 2, 0, 1, 1, 0)
sync_reset;
check_mem(250,"000001001","000110000",2,'1'); -- (0, 0, 0, 2, 2, 1, 0, 0, 1)
sync_reset;
check_mem(251,"000001010","000110000",8,'1'); -- (0, 0, 0, 2, 2, 1, 0, 1, 0)
sync_reset;
check_mem(252,"000001011","000110000",0,'1'); -- (0, 0, 0, 2, 2, 1, 0, 1, 1)
sync_reset;
check_mem(253,"000001100","000110000",8,'1'); -- (0, 0, 0, 2, 2, 1, 1, 0, 0)
sync_reset;
check_mem(254,"000001101","000110000",0,'1'); -- (0, 0, 0, 2, 2, 1, 1, 0, 1)
sync_reset;
check_mem(255,"000001110","000110000",8,'1'); -- (0, 0, 0, 2, 2, 1, 1, 1, 0)
sync_reset;
check_mem(256,"000001110","000110001",0,'1'); -- (0, 0, 0, 2, 2, 1, 1, 1, 2)
sync_reset;
check_mem(257,"000001101","000110010",2,'1'); -- (0, 0, 0, 2, 2, 1, 1, 2, 1)
sync_reset;
check_mem(258,"000001011","000110100",2,'1'); -- (0, 0, 0, 2, 2, 1, 2, 1, 1)
sync_reset;
check_mem(259,"001000000","000000000",4,'1'); -- (0, 0, 1, 0, 0, 0, 0, 0, 0)
sync_reset;
check_mem(260,"001000000","000000001",0,'1'); -- (0, 0, 1, 0, 0, 0, 0, 0, 2)
sync_reset;
check_mem(261,"001000010","000000001",1,'1'); -- (0, 0, 1, 0, 0, 0, 0, 1, 2)
sync_reset;
check_mem(262,"001000000","000000010",0,'1'); -- (0, 0, 1, 0, 0, 0, 0, 2, 0)
sync_reset;
check_mem(263,"001000001","000000010",0,'1'); -- (0, 0, 1, 0, 0, 0, 0, 2, 1)
sync_reset;
check_mem(264,"001000100","000000001",0,'1'); -- (0, 0, 1, 0, 0, 0, 1, 0, 2)
sync_reset;
check_mem(265,"001000100","000000010",4,'1'); -- (0, 0, 1, 0, 0, 0, 1, 2, 0)
sync_reset;
check_mem(266,"001000100","000000011",0,'1'); -- (0, 0, 1, 0, 0, 0, 1, 2, 2)
sync_reset;
check_mem(267,"001000000","000000100",0,'1'); -- (0, 0, 1, 0, 0, 0, 2, 0, 0)
sync_reset;
check_mem(268,"001000001","000000100",0,'1'); -- (0, 0, 1, 0, 0, 0, 2, 0, 1)
sync_reset;
check_mem(269,"001000010","000000100",0,'1'); -- (0, 0, 1, 0, 0, 0, 2, 1, 0)
sync_reset;
check_mem(270,"001000010","000000101",1,'1'); -- (0, 0, 1, 0, 0, 0, 2, 1, 2)
sync_reset;
check_mem(271,"001000001","000000110",0,'1'); -- (0, 0, 1, 0, 0, 0, 2, 2, 1)
sync_reset;
check_mem(272,"001001000","000000001",6,'1'); -- (0, 0, 1, 0, 0, 1, 0, 0, 2)
sync_reset;
check_mem(273,"001001000","000000010",8,'1'); -- (0, 0, 1, 0, 0, 1, 0, 2, 0)
sync_reset;
check_mem(274,"001001000","000000011",0,'1'); -- (0, 0, 1, 0, 0, 1, 0, 2, 2)
sync_reset;
check_mem(275,"001001100","000000011",4,'1'); -- (0, 0, 1, 0, 0, 1, 1, 2, 2)
sync_reset;
check_mem(276,"001001000","000000100",8,'1'); -- (0, 0, 1, 0, 0, 1, 2, 0, 0)
sync_reset;
check_mem(277,"001001000","000000101",0,'1'); -- (0, 0, 1, 0, 0, 1, 2, 0, 2)
sync_reset;
check_mem(278,"001001010","000000101",0,'1'); -- (0, 0, 1, 0, 0, 1, 2, 1, 2)
sync_reset;
check_mem(279,"001001000","000000110",8,'1'); -- (0, 0, 1, 0, 0, 1, 2, 2, 0)
sync_reset;
check_mem(280,"001000000","000001000",0,'1'); -- (0, 0, 1, 0, 0, 2, 0, 0, 0)
sync_reset;
check_mem(281,"001000001","000001000",4,'1'); -- (0, 0, 1, 0, 0, 2, 0, 0, 1)
sync_reset;
check_mem(282,"001000010","000001000",4,'1'); -- (0, 0, 1, 0, 0, 2, 0, 1, 0)
sync_reset;
check_mem(283,"001000010","000001001",0,'1'); -- (0, 0, 1, 0, 0, 2, 0, 1, 2)
sync_reset;
check_mem(284,"001000001","000001010",0,'1'); -- (0, 0, 1, 0, 0, 2, 0, 2, 1)
sync_reset;
check_mem(285,"001000100","000001000",4,'1'); -- (0, 0, 1, 0, 0, 2, 1, 0, 0)
sync_reset;
check_mem(286,"001000100","000001001",0,'1'); -- (0, 0, 1, 0, 0, 2, 1, 0, 2)
sync_reset;
check_mem(287,"001000110","000001001",4,'1'); -- (0, 0, 1, 0, 0, 2, 1, 1, 2)
sync_reset;
check_mem(288,"001000100","000001010",0,'1'); -- (0, 0, 1, 0, 0, 2, 1, 2, 0)
sync_reset;
check_mem(289,"001000101","000001010",4,'1'); -- (0, 0, 1, 0, 0, 2, 1, 2, 1)
sync_reset;
check_mem(290,"001000001","000001100",0,'1'); -- (0, 0, 1, 0, 0, 2, 2, 0, 1)
sync_reset;
check_mem(291,"001000010","000001100",1,'1'); -- (0, 0, 1, 0, 0, 2, 2, 1, 0)
sync_reset;
check_mem(292,"001000011","000001100",3,'1'); -- (0, 0, 1, 0, 0, 2, 2, 1, 1)
sync_reset;
check_mem(293,"001010000","000000001",6,'1'); -- (0, 0, 1, 0, 1, 0, 0, 0, 2)
sync_reset;
check_mem(294,"001010000","000000010",0,'1'); -- (0, 0, 1, 0, 1, 0, 0, 2, 0)
sync_reset;
check_mem(295,"001010000","000000011",6,'1'); -- (0, 0, 1, 0, 1, 0, 0, 2, 2)
sync_reset;
check_mem(296,"001010000","000000100",0,'1'); -- (0, 0, 1, 0, 1, 0, 2, 0, 0)
sync_reset;
check_mem(297,"001010000","000000101",7,'1'); -- (0, 0, 1, 0, 1, 0, 2, 0, 2)
sync_reset;
check_mem(298,"001010010","000000101",1,'1'); -- (0, 0, 1, 0, 1, 0, 2, 1, 2)
sync_reset;
check_mem(299,"001010000","000000110",8,'1'); -- (0, 0, 1, 0, 1, 0, 2, 2, 0)
sync_reset;
check_mem(300,"001010001","000000110",0,'1'); -- (0, 0, 1, 0, 1, 0, 2, 2, 1)
sync_reset;
check_mem(301,"001011000","000000011",6,'1'); -- (0, 0, 1, 0, 1, 1, 0, 2, 2)
sync_reset;
check_mem(302,"001011000","000000101",3,'1'); -- (0, 0, 1, 0, 1, 1, 2, 0, 2)
sync_reset;
check_mem(303,"001011000","000000110",8,'1'); -- (0, 0, 1, 0, 1, 1, 2, 2, 0)
sync_reset;
check_mem(304,"001010000","000001000",0,'1'); -- (0, 0, 1, 0, 1, 2, 0, 0, 0)
sync_reset;
check_mem(305,"001010000","000001001",0,'1'); -- (0, 0, 1, 0, 1, 2, 0, 0, 2)
sync_reset;
check_mem(306,"001010010","000001001",0,'1'); -- (0, 0, 1, 0, 1, 2, 0, 1, 2)
sync_reset;
check_mem(307,"001010000","000001010",0,'1'); -- (0, 0, 1, 0, 1, 2, 0, 2, 0)
sync_reset;
check_mem(308,"001010001","000001010",0,'1'); -- (0, 0, 1, 0, 1, 2, 0, 2, 1)
sync_reset;
check_mem(309,"001010000","000001100",0,'1'); -- (0, 0, 1, 0, 1, 2, 2, 0, 0)
sync_reset;
check_mem(310,"001010001","000001100",0,'1'); -- (0, 0, 1, 0, 1, 2, 2, 0, 1)
sync_reset;
check_mem(311,"001010010","000001100",1,'1'); -- (0, 0, 1, 0, 1, 2, 2, 1, 0)
sync_reset;
check_mem(312,"001010010","000001101",1,'1'); -- (0, 0, 1, 0, 1, 2, 2, 1, 2)
sync_reset;
check_mem(313,"001010001","000001110",0,'1'); -- (0, 0, 1, 0, 1, 2, 2, 2, 1)
sync_reset;
check_mem(314,"001000000","000010000",0,'1'); -- (0, 0, 1, 0, 2, 0, 0, 0, 0)
sync_reset;
check_mem(315,"001000001","000010000",5,'1'); -- (0, 0, 1, 0, 2, 0, 0, 0, 1)
sync_reset;
check_mem(316,"001000010","000010000",3,'1'); -- (0, 0, 1, 0, 2, 0, 0, 1, 0)
sync_reset;
check_mem(317,"001000010","000010001",0,'1'); -- (0, 0, 1, 0, 2, 0, 0, 1, 2)
sync_reset;
check_mem(318,"001000001","000010010",1,'1'); -- (0, 0, 1, 0, 2, 0, 0, 2, 1)
sync_reset;
check_mem(319,"001000100","000010000",1,'1'); -- (0, 0, 1, 0, 2, 0, 1, 0, 0)
sync_reset;
check_mem(320,"001000100","000010001",0,'1'); -- (0, 0, 1, 0, 2, 0, 1, 0, 2)
sync_reset;
check_mem(321,"001000110","000010001",0,'1'); -- (0, 0, 1, 0, 2, 0, 1, 1, 2)
sync_reset;
check_mem(322,"001000100","000010010",1,'1'); -- (0, 0, 1, 0, 2, 0, 1, 2, 0)
sync_reset;
check_mem(323,"001000101","000010010",1,'1'); -- (0, 0, 1, 0, 2, 0, 1, 2, 1)
sync_reset;
check_mem(324,"001000001","000010100",0,'1'); -- (0, 0, 1, 0, 2, 0, 2, 0, 1)
sync_reset;
check_mem(325,"001000010","000010100",0,'1'); -- (0, 0, 1, 0, 2, 0, 2, 1, 0)
sync_reset;
check_mem(326,"001000011","000010100",5,'1'); -- (0, 0, 1, 0, 2, 0, 2, 1, 1)
sync_reset;
check_mem(327,"001001000","000010000",8,'1'); -- (0, 0, 1, 0, 2, 1, 0, 0, 0)
sync_reset;
check_mem(328,"001001000","000010001",0,'1'); -- (0, 0, 1, 0, 2, 1, 0, 0, 2)
sync_reset;
check_mem(329,"001001010","000010001",0,'1'); -- (0, 0, 1, 0, 2, 1, 0, 1, 2)
sync_reset;
check_mem(330,"001001000","000010010",1,'1'); -- (0, 0, 1, 0, 2, 1, 0, 2, 0)
sync_reset;
check_mem(331,"001001100","000010001",0,'1'); -- (0, 0, 1, 0, 2, 1, 1, 0, 2)
sync_reset;
check_mem(332,"001001100","000010010",1,'1'); -- (0, 0, 1, 0, 2, 1, 1, 2, 0)
sync_reset;
check_mem(333,"001001100","000010011",0,'1'); -- (0, 0, 1, 0, 2, 1, 1, 2, 2)
sync_reset;
check_mem(334,"001001000","000010100",0,'1'); -- (0, 0, 1, 0, 2, 1, 2, 0, 0)
sync_reset;
check_mem(335,"001001010","000010100",8,'1'); -- (0, 0, 1, 0, 2, 1, 2, 1, 0)
sync_reset;
check_mem(336,"001001010","000010101",0,'1'); -- (0, 0, 1, 0, 2, 1, 2, 1, 2)
sync_reset;
check_mem(337,"001000001","000011000",3,'1'); -- (0, 0, 1, 0, 2, 2, 0, 0, 1)
sync_reset;
check_mem(338,"001000010","000011000",3,'1'); -- (0, 0, 1, 0, 2, 2, 0, 1, 0)
sync_reset;
check_mem(339,"001000011","000011000",3,'1'); -- (0, 0, 1, 0, 2, 2, 0, 1, 1)
sync_reset;
check_mem(340,"001000100","000011000",3,'1'); -- (0, 0, 1, 0, 2, 2, 1, 0, 0)
sync_reset;
check_mem(341,"001000101","000011000",3,'1'); -- (0, 0, 1, 0, 2, 2, 1, 0, 1)
sync_reset;
check_mem(342,"001000110","000011000",3,'1'); -- (0, 0, 1, 0, 2, 2, 1, 1, 0)
sync_reset;
check_mem(343,"001000110","000011001",0,'1'); -- (0, 0, 1, 0, 2, 2, 1, 1, 2)
sync_reset;
check_mem(344,"001000101","000011010",0,'1'); -- (0, 0, 1, 0, 2, 2, 1, 2, 1)
sync_reset;
check_mem(345,"001000011","000011100",3,'1'); -- (0, 0, 1, 0, 2, 2, 2, 1, 1)
sync_reset;
check_mem(346,"001100000","000000001",6,'1'); -- (0, 0, 1, 1, 0, 0, 0, 0, 2)
sync_reset;
check_mem(347,"001100000","000000010",4,'1'); -- (0, 0, 1, 1, 0, 0, 0, 2, 0)
sync_reset;
check_mem(348,"001100000","000000011",6,'1'); -- (0, 0, 1, 1, 0, 0, 0, 2, 2)
sync_reset;
check_mem(349,"001100100","000000011",0,'1'); -- (0, 0, 1, 1, 0, 0, 1, 2, 2)
sync_reset;
check_mem(350,"001100000","000000100",4,'1'); -- (0, 0, 1, 1, 0, 0, 2, 0, 0)
sync_reset;
check_mem(351,"001100000","000000101",7,'1'); -- (0, 0, 1, 1, 0, 0, 2, 0, 2)
sync_reset;
check_mem(352,"001100010","000000101",1,'1'); -- (0, 0, 1, 1, 0, 0, 2, 1, 2)
sync_reset;
check_mem(353,"001100000","000000110",8,'1'); -- (0, 0, 1, 1, 0, 0, 2, 2, 0)
sync_reset;
check_mem(354,"001100001","000000110",0,'1'); -- (0, 0, 1, 1, 0, 0, 2, 2, 1)
sync_reset;
check_mem(355,"001101000","000000011",4,'1'); -- (0, 0, 1, 1, 0, 1, 0, 2, 2)
sync_reset;
check_mem(356,"001101000","000000101",4,'1'); -- (0, 0, 1, 1, 0, 1, 2, 0, 2)
sync_reset;
check_mem(357,"001101000","000000110",8,'1'); -- (0, 0, 1, 1, 0, 1, 2, 2, 0)
sync_reset;
check_mem(358,"001100000","000001000",0,'1'); -- (0, 0, 1, 1, 0, 2, 0, 0, 0)
sync_reset;
check_mem(359,"001100000","000001001",0,'1'); -- (0, 0, 1, 1, 0, 2, 0, 0, 2)
sync_reset;
check_mem(360,"001100010","000001001",0,'1'); -- (0, 0, 1, 1, 0, 2, 0, 1, 2)
sync_reset;
check_mem(361,"001100000","000001010",0,'1'); -- (0, 0, 1, 1, 0, 2, 0, 2, 0)
sync_reset;
check_mem(362,"001100001","000001010",0,'1'); -- (0, 0, 1, 1, 0, 2, 0, 2, 1)
sync_reset;
check_mem(363,"001100100","000001001",0,'1'); -- (0, 0, 1, 1, 0, 2, 1, 0, 2)
sync_reset;
check_mem(364,"001100100","000001010",0,'1'); -- (0, 0, 1, 1, 0, 2, 1, 2, 0)
sync_reset;
check_mem(365,"001100100","000001011",0,'1'); -- (0, 0, 1, 1, 0, 2, 1, 2, 2)
sync_reset;
check_mem(366,"001100000","000001100",0,'1'); -- (0, 0, 1, 1, 0, 2, 2, 0, 0)
sync_reset;
check_mem(367,"001100001","000001100",0,'1'); -- (0, 0, 1, 1, 0, 2, 2, 0, 1)
sync_reset;
check_mem(368,"001100010","000001100",0,'1'); -- (0, 0, 1, 1, 0, 2, 2, 1, 0)
sync_reset;
check_mem(369,"001100010","000001101",1,'1'); -- (0, 0, 1, 1, 0, 2, 2, 1, 2)
sync_reset;
check_mem(370,"001100001","000001110",0,'1'); -- (0, 0, 1, 1, 0, 2, 2, 2, 1)
sync_reset;
check_mem(371,"001110000","000000011",6,'1'); -- (0, 0, 1, 1, 1, 0, 0, 2, 2)
sync_reset;
check_mem(372,"001110000","000000101",7,'1'); -- (0, 0, 1, 1, 1, 0, 2, 0, 2)
sync_reset;
check_mem(373,"001110000","000000110",8,'1'); -- (0, 0, 1, 1, 1, 0, 2, 2, 0)
sync_reset;
check_mem(374,"001110000","000001001",6,'1'); -- (0, 0, 1, 1, 1, 2, 0, 0, 2)
sync_reset;
check_mem(375,"001110000","000001010",6,'1'); -- (0, 0, 1, 1, 1, 2, 0, 2, 0)
sync_reset;
check_mem(376,"001110000","000001011",6,'1'); -- (0, 0, 1, 1, 1, 2, 0, 2, 2)
sync_reset;
check_mem(377,"001110000","000001100",0,'1'); -- (0, 0, 1, 1, 1, 2, 2, 0, 0)
sync_reset;
check_mem(378,"001110000","000001101",7,'1'); -- (0, 0, 1, 1, 1, 2, 2, 0, 2)
sync_reset;
check_mem(379,"001110010","000001101",1,'1'); -- (0, 0, 1, 1, 1, 2, 2, 1, 2)
sync_reset;
check_mem(380,"001110000","000001110",8,'1'); -- (0, 0, 1, 1, 1, 2, 2, 2, 0)
sync_reset;
check_mem(381,"001110001","000001110",0,'1'); -- (0, 0, 1, 1, 1, 2, 2, 2, 1)
sync_reset;
check_mem(382,"001100000","000010000",0,'1'); -- (0, 0, 1, 1, 2, 0, 0, 0, 0)
sync_reset;
check_mem(383,"001100000","000010001",0,'1'); -- (0, 0, 1, 1, 2, 0, 0, 0, 2)
sync_reset;
check_mem(384,"001100010","000010001",0,'1'); -- (0, 0, 1, 1, 2, 0, 0, 1, 2)
sync_reset;
check_mem(385,"001100000","000010010",1,'1'); -- (0, 0, 1, 1, 2, 0, 0, 2, 0)
sync_reset;
check_mem(386,"001100001","000010010",1,'1'); -- (0, 0, 1, 1, 2, 0, 0, 2, 1)
sync_reset;
check_mem(387,"001100100","000010001",0,'1'); -- (0, 0, 1, 1, 2, 0, 1, 0, 2)
sync_reset;
check_mem(388,"001100100","000010010",0,'1'); -- (0, 0, 1, 1, 2, 0, 1, 2, 0)
sync_reset;
check_mem(389,"001100100","000010011",0,'1'); -- (0, 0, 1, 1, 2, 0, 1, 2, 2)
sync_reset;
check_mem(390,"001100000","000010100",0,'1'); -- (0, 0, 1, 1, 2, 0, 2, 0, 0)
sync_reset;
check_mem(391,"001100001","000010100",5,'1'); -- (0, 0, 1, 1, 2, 0, 2, 0, 1)
sync_reset;
check_mem(392,"001100010","000010100",0,'1'); -- (0, 0, 1, 1, 2, 0, 2, 1, 0)
sync_reset;
check_mem(393,"001100010","000010101",0,'1'); -- (0, 0, 1, 1, 2, 0, 2, 1, 2)
sync_reset;
check_mem(394,"001100001","000010110",1,'1'); -- (0, 0, 1, 1, 2, 0, 2, 2, 1)
sync_reset;
check_mem(395,"001101000","000010001",0,'1'); -- (0, 0, 1, 1, 2, 1, 0, 0, 2)
sync_reset;
check_mem(396,"001101000","000010010",1,'1'); -- (0, 0, 1, 1, 2, 1, 0, 2, 0)
sync_reset;
check_mem(397,"001101000","000010011",0,'1'); -- (0, 0, 1, 1, 2, 1, 0, 2, 2)
sync_reset;
check_mem(398,"001101100","000010011",0,'1'); -- (0, 0, 1, 1, 2, 1, 1, 2, 2)
sync_reset;
check_mem(399,"001101000","000010100",8,'1'); -- (0, 0, 1, 1, 2, 1, 2, 0, 0)
sync_reset;
check_mem(400,"001101000","000010101",0,'1'); -- (0, 0, 1, 1, 2, 1, 2, 0, 2)
sync_reset;
check_mem(401,"001101010","000010101",0,'1'); -- (0, 0, 1, 1, 2, 1, 2, 1, 2)
sync_reset;
check_mem(402,"001101000","000010110",8,'1'); -- (0, 0, 1, 1, 2, 1, 2, 2, 0)
sync_reset;
check_mem(403,"001100000","000011000",0,'1'); -- (0, 0, 1, 1, 2, 2, 0, 0, 0)
sync_reset;
check_mem(404,"001100001","000011000",0,'1'); -- (0, 0, 1, 1, 2, 2, 0, 0, 1)
sync_reset;
check_mem(405,"001100010","000011000",0,'1'); -- (0, 0, 1, 1, 2, 2, 0, 1, 0)
sync_reset;
check_mem(406,"001100010","000011001",0,'1'); -- (0, 0, 1, 1, 2, 2, 0, 1, 2)
sync_reset;
check_mem(407,"001100001","000011010",1,'1'); -- (0, 0, 1, 1, 2, 2, 0, 2, 1)
sync_reset;
check_mem(408,"001100100","000011000",0,'1'); -- (0, 0, 1, 1, 2, 2, 1, 0, 0)
sync_reset;
check_mem(409,"001100100","000011001",0,'1'); -- (0, 0, 1, 1, 2, 2, 1, 0, 2)
sync_reset;
check_mem(410,"001100110","000011001",0,'1'); -- (0, 0, 1, 1, 2, 2, 1, 1, 2)
sync_reset;
check_mem(411,"001100100","000011010",0,'1'); -- (0, 0, 1, 1, 2, 2, 1, 2, 0)
sync_reset;
check_mem(412,"001100101","000011010",1,'1'); -- (0, 0, 1, 1, 2, 2, 1, 2, 1)
sync_reset;
check_mem(413,"001100001","000011100",0,'1'); -- (0, 0, 1, 1, 2, 2, 2, 0, 1)
sync_reset;
check_mem(414,"001100010","000011100",0,'1'); -- (0, 0, 1, 1, 2, 2, 2, 1, 0)
sync_reset;
check_mem(415,"001100011","000011100",0,'1'); -- (0, 0, 1, 1, 2, 2, 2, 1, 1)
sync_reset;
check_mem(416,"001000000","000100000",0,'1'); -- (0, 0, 1, 2, 0, 0, 0, 0, 0)
sync_reset;
check_mem(417,"001000001","000100000",0,'1'); -- (0, 0, 1, 2, 0, 0, 0, 0, 1)
sync_reset;
check_mem(418,"001000010","000100000",4,'1'); -- (0, 0, 1, 2, 0, 0, 0, 1, 0)
sync_reset;
check_mem(419,"001000010","000100001",1,'1'); -- (0, 0, 1, 2, 0, 0, 0, 1, 2)
sync_reset;
check_mem(420,"001000001","000100010",0,'1'); -- (0, 0, 1, 2, 0, 0, 0, 2, 1)
sync_reset;
check_mem(421,"001000100","000100000",4,'1'); -- (0, 0, 1, 2, 0, 0, 1, 0, 0)
sync_reset;
check_mem(422,"001000100","000100001",0,'1'); -- (0, 0, 1, 2, 0, 0, 1, 0, 2)
sync_reset;
check_mem(423,"001000110","000100001",4,'1'); -- (0, 0, 1, 2, 0, 0, 1, 1, 2)
sync_reset;
check_mem(424,"001000100","000100010",0,'1'); -- (0, 0, 1, 2, 0, 0, 1, 2, 0)
sync_reset;
check_mem(425,"001000101","000100010",0,'1'); -- (0, 0, 1, 2, 0, 0, 1, 2, 1)
sync_reset;
check_mem(426,"001000001","000100100",0,'1'); -- (0, 0, 1, 2, 0, 0, 2, 0, 1)
sync_reset;
check_mem(427,"001000010","000100100",0,'1'); -- (0, 0, 1, 2, 0, 0, 2, 1, 0)
sync_reset;
check_mem(428,"001000011","000100100",0,'1'); -- (0, 0, 1, 2, 0, 0, 2, 1, 1)
sync_reset;
check_mem(429,"001001000","000100000",8,'1'); -- (0, 0, 1, 2, 0, 1, 0, 0, 0)
sync_reset;
check_mem(430,"001001000","000100001",0,'1'); -- (0, 0, 1, 2, 0, 1, 0, 0, 2)
sync_reset;
check_mem(431,"001001010","000100001",0,'1'); -- (0, 0, 1, 2, 0, 1, 0, 1, 2)
sync_reset;
check_mem(432,"001001000","000100010",0,'1'); -- (0, 0, 1, 2, 0, 1, 0, 2, 0)
sync_reset;
check_mem(433,"001001100","000100001",4,'1'); -- (0, 0, 1, 2, 0, 1, 1, 0, 2)
sync_reset;
check_mem(434,"001001100","000100010",0,'1'); -- (0, 0, 1, 2, 0, 1, 1, 2, 0)
sync_reset;
check_mem(435,"001001100","000100011",0,'1'); -- (0, 0, 1, 2, 0, 1, 1, 2, 2)
sync_reset;
check_mem(436,"001001000","000100100",0,'1'); -- (0, 0, 1, 2, 0, 1, 2, 0, 0)
sync_reset;
check_mem(437,"001001010","000100100",0,'1'); -- (0, 0, 1, 2, 0, 1, 2, 1, 0)
sync_reset;
check_mem(438,"001001010","000100101",0,'1'); -- (0, 0, 1, 2, 0, 1, 2, 1, 2)
sync_reset;
check_mem(439,"001000001","000101000",4,'1'); -- (0, 0, 1, 2, 0, 2, 0, 0, 1)
sync_reset;
check_mem(440,"001000010","000101000",4,'1'); -- (0, 0, 1, 2, 0, 2, 0, 1, 0)
sync_reset;
check_mem(441,"001000011","000101000",4,'1'); -- (0, 0, 1, 2, 0, 2, 0, 1, 1)
sync_reset;
check_mem(442,"001000100","000101000",4,'1'); -- (0, 0, 1, 2, 0, 2, 1, 0, 0)
sync_reset;
check_mem(443,"001000101","000101000",4,'1'); -- (0, 0, 1, 2, 0, 2, 1, 0, 1)
sync_reset;
check_mem(444,"001000110","000101000",4,'1'); -- (0, 0, 1, 2, 0, 2, 1, 1, 0)
sync_reset;
check_mem(445,"001000110","000101001",4,'1'); -- (0, 0, 1, 2, 0, 2, 1, 1, 2)
sync_reset;
check_mem(446,"001000101","000101010",4,'1'); -- (0, 0, 1, 2, 0, 2, 1, 2, 1)
sync_reset;
check_mem(447,"001000011","000101100",0,'1'); -- (0, 0, 1, 2, 0, 2, 2, 1, 1)
sync_reset;
check_mem(448,"001010000","000100000",0,'1'); -- (0, 0, 1, 2, 1, 0, 0, 0, 0)
sync_reset;
check_mem(449,"001010000","000100001",0,'1'); -- (0, 0, 1, 2, 1, 0, 0, 0, 2)
sync_reset;
check_mem(450,"001010010","000100001",0,'1'); -- (0, 0, 1, 2, 1, 0, 0, 1, 2)
sync_reset;
check_mem(451,"001010000","000100010",0,'1'); -- (0, 0, 1, 2, 1, 0, 0, 2, 0)
sync_reset;
check_mem(452,"001010001","000100010",0,'1'); -- (0, 0, 1, 2, 1, 0, 0, 2, 1)
sync_reset;
check_mem(453,"001010000","000100100",0,'1'); -- (0, 0, 1, 2, 1, 0, 2, 0, 0)
sync_reset;
check_mem(454,"001010001","000100100",0,'1'); -- (0, 0, 1, 2, 1, 0, 2, 0, 1)
sync_reset;
check_mem(455,"001010010","000100100",0,'1'); -- (0, 0, 1, 2, 1, 0, 2, 1, 0)
sync_reset;
check_mem(456,"001010010","000100101",1,'1'); -- (0, 0, 1, 2, 1, 0, 2, 1, 2)
sync_reset;
check_mem(457,"001010001","000100110",0,'1'); -- (0, 0, 1, 2, 1, 0, 2, 2, 1)
sync_reset;
check_mem(458,"001011000","000100001",6,'1'); -- (0, 0, 1, 2, 1, 1, 0, 0, 2)
sync_reset;
check_mem(459,"001011000","000100010",0,'1'); -- (0, 0, 1, 2, 1, 1, 0, 2, 0)
sync_reset;
check_mem(460,"001011000","000100011",6,'1'); -- (0, 0, 1, 2, 1, 1, 0, 2, 2)
sync_reset;
check_mem(461,"001011000","000100100",0,'1'); -- (0, 0, 1, 2, 1, 1, 2, 0, 0)
sync_reset;
check_mem(462,"001011000","000100101",0,'1'); -- (0, 0, 1, 2, 1, 1, 2, 0, 2)
sync_reset;
check_mem(463,"001011010","000100101",0,'1'); -- (0, 0, 1, 2, 1, 1, 2, 1, 2)
sync_reset;
check_mem(464,"001011000","000100110",8,'1'); -- (0, 0, 1, 2, 1, 1, 2, 2, 0)
sync_reset;
check_mem(465,"001010000","000101000",0,'1'); -- (0, 0, 1, 2, 1, 2, 0, 0, 0)
sync_reset;
check_mem(466,"001010001","000101000",0,'1'); -- (0, 0, 1, 2, 1, 2, 0, 0, 1)
sync_reset;
check_mem(467,"001010010","000101000",0,'1'); -- (0, 0, 1, 2, 1, 2, 0, 1, 0)
sync_reset;
check_mem(468,"001010010","000101001",0,'1'); -- (0, 0, 1, 2, 1, 2, 0, 1, 2)
sync_reset;
check_mem(469,"001010001","000101010",0,'1'); -- (0, 0, 1, 2, 1, 2, 0, 2, 1)
sync_reset;
check_mem(470,"001010001","000101100",0,'1'); -- (0, 0, 1, 2, 1, 2, 2, 0, 1)
sync_reset;
check_mem(471,"001010010","000101100",0,'1'); -- (0, 0, 1, 2, 1, 2, 2, 1, 0)
sync_reset;
check_mem(472,"001010011","000101100",0,'1'); -- (0, 0, 1, 2, 1, 2, 2, 1, 1)
sync_reset;
check_mem(473,"001000001","000110000",5,'1'); -- (0, 0, 1, 2, 2, 0, 0, 0, 1)
sync_reset;
check_mem(474,"001000010","000110000",5,'1'); -- (0, 0, 1, 2, 2, 0, 0, 1, 0)
sync_reset;
check_mem(475,"001000011","000110000",5,'1'); -- (0, 0, 1, 2, 2, 0, 0, 1, 1)
sync_reset;
check_mem(476,"001000100","000110000",5,'1'); -- (0, 0, 1, 2, 2, 0, 1, 0, 0)
sync_reset;
check_mem(477,"001000101","000110000",5,'1'); -- (0, 0, 1, 2, 2, 0, 1, 0, 1)
sync_reset;
check_mem(478,"001000110","000110000",5,'1'); -- (0, 0, 1, 2, 2, 0, 1, 1, 0)
sync_reset;
check_mem(479,"001000110","000110001",0,'1'); -- (0, 0, 1, 2, 2, 0, 1, 1, 2)
sync_reset;
check_mem(480,"001000101","000110010",5,'1'); -- (0, 0, 1, 2, 2, 0, 1, 2, 1)
sync_reset;
check_mem(481,"001000011","000110100",5,'1'); -- (0, 0, 1, 2, 2, 0, 2, 1, 1)
sync_reset;
check_mem(482,"001001000","000110000",0,'1'); -- (0, 0, 1, 2, 2, 1, 0, 0, 0)
sync_reset;
check_mem(483,"001001010","000110000",8,'1'); -- (0, 0, 1, 2, 2, 1, 0, 1, 0)
sync_reset;
check_mem(484,"001001010","000110001",0,'1'); -- (0, 0, 1, 2, 2, 1, 0, 1, 2)
sync_reset;
check_mem(485,"001001100","000110000",8,'1'); -- (0, 0, 1, 2, 2, 1, 1, 0, 0)
sync_reset;
check_mem(486,"001001100","000110001",0,'1'); -- (0, 0, 1, 2, 2, 1, 1, 0, 2)
sync_reset;
check_mem(487,"001001110","000110001",0,'1'); -- (0, 0, 1, 2, 2, 1, 1, 1, 2)
sync_reset;
check_mem(488,"001001100","000110010",1,'1'); -- (0, 0, 1, 2, 2, 1, 1, 2, 0)
sync_reset;
check_mem(489,"001001010","000110100",0,'1'); -- (0, 0, 1, 2, 2, 1, 2, 1, 0)
sync_reset;
check_mem(490,"000000001","001000000",0,'1'); -- (0, 0, 2, 0, 0, 0, 0, 0, 1)
sync_reset;
check_mem(491,"000000010","001000000",8,'1'); -- (0, 0, 2, 0, 0, 0, 0, 1, 0)
sync_reset;
check_mem(492,"000000011","001000000",0,'1'); -- (0, 0, 2, 0, 0, 0, 0, 1, 1)
sync_reset;
check_mem(493,"000000100","001000000",0,'1'); -- (0, 0, 2, 0, 0, 0, 1, 0, 0)
sync_reset;
check_mem(494,"000000101","001000000",0,'1'); -- (0, 0, 2, 0, 0, 0, 1, 0, 1)
sync_reset;
check_mem(495,"000000110","001000000",8,'1'); -- (0, 0, 2, 0, 0, 0, 1, 1, 0)
sync_reset;
check_mem(496,"000000110","001000001",0,'1'); -- (0, 0, 2, 0, 0, 0, 1, 1, 2)
sync_reset;
check_mem(497,"000000101","001000010",0,'1'); -- (0, 0, 2, 0, 0, 0, 1, 2, 1)
sync_reset;
check_mem(498,"000000011","001000100",4,'1'); -- (0, 0, 2, 0, 0, 0, 2, 1, 1)
sync_reset;
check_mem(499,"000001000","001000000",0,'1'); -- (0, 0, 2, 0, 0, 1, 0, 0, 0)
sync_reset;
check_mem(500,"000001001","001000000",0,'1'); -- (0, 0, 2, 0, 0, 1, 0, 0, 1)
sync_reset;
check_mem(501,"000001010","001000000",0,'1'); -- (0, 0, 2, 0, 0, 1, 0, 1, 0)
sync_reset;
check_mem(502,"000001010","001000001",4,'1'); -- (0, 0, 2, 0, 0, 1, 0, 1, 2)
sync_reset;
check_mem(503,"000001001","001000010",4,'1'); -- (0, 0, 2, 0, 0, 1, 0, 2, 1)
sync_reset;
check_mem(504,"000001100","001000000",0,'1'); -- (0, 0, 2, 0, 0, 1, 1, 0, 0)
sync_reset;
check_mem(505,"000001100","001000001",3,'1'); -- (0, 0, 2, 0, 0, 1, 1, 0, 2)
sync_reset;
check_mem(506,"000001110","001000001",0,'1'); -- (0, 0, 2, 0, 0, 1, 1, 1, 2)
sync_reset;
check_mem(507,"000001100","001000010",3,'1'); -- (0, 0, 2, 0, 0, 1, 1, 2, 0)
sync_reset;
check_mem(508,"000001101","001000010",1,'1'); -- (0, 0, 2, 0, 0, 1, 1, 2, 1)
sync_reset;
check_mem(509,"000001001","001000100",4,'1'); -- (0, 0, 2, 0, 0, 1, 2, 0, 1)
sync_reset;
check_mem(510,"000001010","001000100",4,'1'); -- (0, 0, 2, 0, 0, 1, 2, 1, 0)
sync_reset;
check_mem(511,"000001011","001000100",0,'1'); -- (0, 0, 2, 0, 0, 1, 2, 1, 1)
sync_reset;
check_mem(512,"000000011","001001000",0,'1'); -- (0, 0, 2, 0, 0, 2, 0, 1, 1)
sync_reset;
check_mem(513,"000000101","001001000",0,'1'); -- (0, 0, 2, 0, 0, 2, 1, 0, 1)
sync_reset;
check_mem(514,"000000110","001001000",8,'1'); -- (0, 0, 2, 0, 0, 2, 1, 1, 0)
sync_reset;
check_mem(515,"000010000","001000000",0,'1'); -- (0, 0, 2, 0, 1, 0, 0, 0, 0)
sync_reset;
check_mem(516,"000010001","001000000",0,'1'); -- (0, 0, 2, 0, 1, 0, 0, 0, 1)
sync_reset;
check_mem(517,"000010010","001000000",1,'1'); -- (0, 0, 2, 0, 1, 0, 0, 1, 0)
sync_reset;
check_mem(518,"000010010","001000001",1,'1'); -- (0, 0, 2, 0, 1, 0, 0, 1, 2)
sync_reset;
check_mem(519,"000010001","001000010",0,'1'); -- (0, 0, 2, 0, 1, 0, 0, 2, 1)
sync_reset;
check_mem(520,"000010100","001000000",0,'1'); -- (0, 0, 2, 0, 1, 0, 1, 0, 0)
sync_reset;
check_mem(521,"000010100","001000001",5,'1'); -- (0, 0, 2, 0, 1, 0, 1, 0, 2)
sync_reset;
check_mem(522,"000010110","001000001",1,'1'); -- (0, 0, 2, 0, 1, 0, 1, 1, 2)
sync_reset;
check_mem(523,"000010100","001000010",0,'1'); -- (0, 0, 2, 0, 1, 0, 1, 2, 0)
sync_reset;
check_mem(524,"000010101","001000010",0,'1'); -- (0, 0, 2, 0, 1, 0, 1, 2, 1)
sync_reset;
check_mem(525,"000010001","001000100",0,'1'); -- (0, 0, 2, 0, 1, 0, 2, 0, 1)
sync_reset;
check_mem(526,"000010010","001000100",0,'1'); -- (0, 0, 2, 0, 1, 0, 2, 1, 0)
sync_reset;
check_mem(527,"000010011","001000100",0,'1'); -- (0, 0, 2, 0, 1, 0, 2, 1, 1)
sync_reset;
check_mem(528,"000011000","001000000",3,'1'); -- (0, 0, 2, 0, 1, 1, 0, 0, 0)
sync_reset;
check_mem(529,"000011000","001000001",1,'1'); -- (0, 0, 2, 0, 1, 1, 0, 0, 2)
sync_reset;
check_mem(530,"000011010","001000001",0,'1'); -- (0, 0, 2, 0, 1, 1, 0, 1, 2)
sync_reset;
check_mem(531,"000011000","001000010",0,'1'); -- (0, 0, 2, 0, 1, 1, 0, 2, 0)
sync_reset;
check_mem(532,"000011001","001000010",0,'1'); -- (0, 0, 2, 0, 1, 1, 0, 2, 1)
sync_reset;
check_mem(533,"000011100","001000001",3,'1'); -- (0, 0, 2, 0, 1, 1, 1, 0, 2)
sync_reset;
check_mem(534,"000011100","001000010",3,'1'); -- (0, 0, 2, 0, 1, 1, 1, 2, 0)
sync_reset;
check_mem(535,"000011100","001000011",3,'1'); -- (0, 0, 2, 0, 1, 1, 1, 2, 2)
sync_reset;
check_mem(536,"000011000","001000100",0,'1'); -- (0, 0, 2, 0, 1, 1, 2, 0, 0)
sync_reset;
check_mem(537,"000011001","001000100",0,'1'); -- (0, 0, 2, 0, 1, 1, 2, 0, 1)
sync_reset;
check_mem(538,"000011010","001000100",0,'1'); -- (0, 0, 2, 0, 1, 1, 2, 1, 0)
sync_reset;
check_mem(539,"000011010","001000101",0,'1'); -- (0, 0, 2, 0, 1, 1, 2, 1, 2)
sync_reset;
check_mem(540,"000011001","001000110",0,'1'); -- (0, 0, 2, 0, 1, 1, 2, 2, 1)
sync_reset;
check_mem(541,"000010001","001001000",0,'1'); -- (0, 0, 2, 0, 1, 2, 0, 0, 1)
sync_reset;
check_mem(542,"000010010","001001000",1,'1'); -- (0, 0, 2, 0, 1, 2, 0, 1, 0)
sync_reset;
check_mem(543,"000010011","001001000",0,'1'); -- (0, 0, 2, 0, 1, 2, 0, 1, 1)
sync_reset;
check_mem(544,"000010100","001001000",8,'1'); -- (0, 0, 2, 0, 1, 2, 1, 0, 0)
sync_reset;
check_mem(545,"000010101","001001000",0,'1'); -- (0, 0, 2, 0, 1, 2, 1, 0, 1)
sync_reset;
check_mem(546,"000010110","001001000",8,'1'); -- (0, 0, 2, 0, 1, 2, 1, 1, 0)
sync_reset;
check_mem(547,"000010101","001001010",0,'1'); -- (0, 0, 2, 0, 1, 2, 1, 2, 1)
sync_reset;
check_mem(548,"000010011","001001100",0,'1'); -- (0, 0, 2, 0, 1, 2, 2, 1, 1)
sync_reset;
check_mem(549,"000000011","001010000",6,'1'); -- (0, 0, 2, 0, 2, 0, 0, 1, 1)
sync_reset;
check_mem(550,"000000101","001010000",0,'1'); -- (0, 0, 2, 0, 2, 0, 1, 0, 1)
sync_reset;
check_mem(551,"000000110","001010000",0,'1'); -- (0, 0, 2, 0, 2, 0, 1, 1, 0)
sync_reset;
check_mem(552,"000001001","001010000",6,'1'); -- (0, 0, 2, 0, 2, 1, 0, 0, 1)
sync_reset;
check_mem(553,"000001010","001010000",6,'1'); -- (0, 0, 2, 0, 2, 1, 0, 1, 0)
sync_reset;
check_mem(554,"000001011","001010000",6,'1'); -- (0, 0, 2, 0, 2, 1, 0, 1, 1)
sync_reset;
check_mem(555,"000001100","001010000",0,'1'); -- (0, 0, 2, 0, 2, 1, 1, 0, 0)
sync_reset;
check_mem(556,"000001101","001010000",7,'1'); -- (0, 0, 2, 0, 2, 1, 1, 0, 1)
sync_reset;
check_mem(557,"000001110","001010000",8,'1'); -- (0, 0, 2, 0, 2, 1, 1, 1, 0)
sync_reset;
check_mem(558,"000001110","001010001",0,'1'); -- (0, 0, 2, 0, 2, 1, 1, 1, 2)
sync_reset;
check_mem(559,"000001101","001010010",1,'1'); -- (0, 0, 2, 0, 2, 1, 1, 2, 1)
sync_reset;
check_mem(560,"000100000","001000000",0,'1'); -- (0, 0, 2, 1, 0, 0, 0, 0, 0)
sync_reset;
check_mem(561,"000100001","001000000",0,'1'); -- (0, 0, 2, 1, 0, 0, 0, 0, 1)
sync_reset;
check_mem(562,"000100010","001000000",0,'1'); -- (0, 0, 2, 1, 0, 0, 0, 1, 0)
sync_reset;
check_mem(563,"000100010","001000001",0,'1'); -- (0, 0, 2, 1, 0, 0, 0, 1, 2)
sync_reset;
check_mem(564,"000100001","001000010",0,'1'); -- (0, 0, 2, 1, 0, 0, 0, 2, 1)
sync_reset;
check_mem(565,"000100100","001000000",0,'1'); -- (0, 0, 2, 1, 0, 0, 1, 0, 0)
sync_reset;
check_mem(566,"000100100","001000001",0,'1'); -- (0, 0, 2, 1, 0, 0, 1, 0, 2)
sync_reset;
check_mem(567,"000100110","001000001",0,'1'); -- (0, 0, 2, 1, 0, 0, 1, 1, 2)
sync_reset;
check_mem(568,"000100100","001000010",0,'1'); -- (0, 0, 2, 1, 0, 0, 1, 2, 0)
sync_reset;
check_mem(569,"000100101","001000010",0,'1'); -- (0, 0, 2, 1, 0, 0, 1, 2, 1)
sync_reset;
check_mem(570,"000100001","001000100",4,'1'); -- (0, 0, 2, 1, 0, 0, 2, 0, 1)
sync_reset;
check_mem(571,"000100010","001000100",4,'1'); -- (0, 0, 2, 1, 0, 0, 2, 1, 0)
sync_reset;
check_mem(572,"000100011","001000100",0,'1'); -- (0, 0, 2, 1, 0, 0, 2, 1, 1)
sync_reset;
check_mem(573,"000101000","001000000",4,'1'); -- (0, 0, 2, 1, 0, 1, 0, 0, 0)
sync_reset;
check_mem(574,"000101000","001000001",0,'1'); -- (0, 0, 2, 1, 0, 1, 0, 0, 2)
sync_reset;
check_mem(575,"000101010","001000001",4,'1'); -- (0, 0, 2, 1, 0, 1, 0, 1, 2)
sync_reset;
check_mem(576,"000101000","001000010",0,'1'); -- (0, 0, 2, 1, 0, 1, 0, 2, 0)
sync_reset;
check_mem(577,"000101001","001000010",4,'1'); -- (0, 0, 2, 1, 0, 1, 0, 2, 1)
sync_reset;
check_mem(578,"000101100","001000001",0,'1'); -- (0, 0, 2, 1, 0, 1, 1, 0, 2)
sync_reset;
check_mem(579,"000101100","001000010",0,'1'); -- (0, 0, 2, 1, 0, 1, 1, 2, 0)
sync_reset;
check_mem(580,"000101100","001000011",0,'1'); -- (0, 0, 2, 1, 0, 1, 1, 2, 2)
sync_reset;
check_mem(581,"000101000","001000100",4,'1'); -- (0, 0, 2, 1, 0, 1, 2, 0, 0)
sync_reset;
check_mem(582,"000101001","001000100",4,'1'); -- (0, 0, 2, 1, 0, 1, 2, 0, 1)
sync_reset;
check_mem(583,"000101010","001000100",4,'1'); -- (0, 0, 2, 1, 0, 1, 2, 1, 0)
sync_reset;
check_mem(584,"000101010","001000101",4,'1'); -- (0, 0, 2, 1, 0, 1, 2, 1, 2)
sync_reset;
check_mem(585,"000101001","001000110",4,'1'); -- (0, 0, 2, 1, 0, 1, 2, 2, 1)
sync_reset;
check_mem(586,"000100001","001001000",0,'1'); -- (0, 0, 2, 1, 0, 2, 0, 0, 1)
sync_reset;
check_mem(587,"000100010","001001000",8,'1'); -- (0, 0, 2, 1, 0, 2, 0, 1, 0)
sync_reset;
check_mem(588,"000100011","001001000",0,'1'); -- (0, 0, 2, 1, 0, 2, 0, 1, 1)
sync_reset;
check_mem(589,"000100100","001001000",0,'1'); -- (0, 0, 2, 1, 0, 2, 1, 0, 0)
sync_reset;
check_mem(590,"000100101","001001000",0,'1'); -- (0, 0, 2, 1, 0, 2, 1, 0, 1)
sync_reset;
check_mem(591,"000100110","001001000",8,'1'); -- (0, 0, 2, 1, 0, 2, 1, 1, 0)
sync_reset;
check_mem(592,"000100101","001001010",0,'1'); -- (0, 0, 2, 1, 0, 2, 1, 2, 1)
sync_reset;
check_mem(593,"000100011","001001100",4,'1'); -- (0, 0, 2, 1, 0, 2, 2, 1, 1)
sync_reset;
check_mem(594,"000110000","001000000",5,'1'); -- (0, 0, 2, 1, 1, 0, 0, 0, 0)
sync_reset;
check_mem(595,"000110000","001000001",5,'1'); -- (0, 0, 2, 1, 1, 0, 0, 0, 2)
sync_reset;
check_mem(596,"000110010","001000001",5,'1'); -- (0, 0, 2, 1, 1, 0, 0, 1, 2)
sync_reset;
check_mem(597,"000110000","001000010",0,'1'); -- (0, 0, 2, 1, 1, 0, 0, 2, 0)
sync_reset;
check_mem(598,"000110001","001000010",0,'1'); -- (0, 0, 2, 1, 1, 0, 0, 2, 1)
sync_reset;
check_mem(599,"000110100","001000001",5,'1'); -- (0, 0, 2, 1, 1, 0, 1, 0, 2)
sync_reset;
check_mem(600,"000110100","001000010",0,'1'); -- (0, 0, 2, 1, 1, 0, 1, 2, 0)
sync_reset;
check_mem(601,"000110100","001000011",0,'1'); -- (0, 0, 2, 1, 1, 0, 1, 2, 2)
sync_reset;
check_mem(602,"000110000","001000100",0,'1'); -- (0, 0, 2, 1, 1, 0, 2, 0, 0)
sync_reset;
check_mem(603,"000110001","001000100",0,'1'); -- (0, 0, 2, 1, 1, 0, 2, 0, 1)
sync_reset;
check_mem(604,"000110010","001000100",0,'1'); -- (0, 0, 2, 1, 1, 0, 2, 1, 0)
sync_reset;
check_mem(605,"000110010","001000101",1,'1'); -- (0, 0, 2, 1, 1, 0, 2, 1, 2)
sync_reset;
check_mem(606,"000110001","001000110",0,'1'); -- (0, 0, 2, 1, 1, 0, 2, 2, 1)
sync_reset;
check_mem(607,"000110000","001001000",8,'1'); -- (0, 0, 2, 1, 1, 2, 0, 0, 0)
sync_reset;
check_mem(608,"000110001","001001000",0,'1'); -- (0, 0, 2, 1, 1, 2, 0, 0, 1)
sync_reset;
check_mem(609,"000110010","001001000",1,'1'); -- (0, 0, 2, 1, 1, 2, 0, 1, 0)
sync_reset;
check_mem(610,"000110001","001001010",0,'1'); -- (0, 0, 2, 1, 1, 2, 0, 2, 1)
sync_reset;
check_mem(611,"000110100","001001000",0,'1'); -- (0, 0, 2, 1, 1, 2, 1, 0, 0)
sync_reset;
check_mem(612,"000110100","001001010",0,'1'); -- (0, 0, 2, 1, 1, 2, 1, 2, 0)
sync_reset;
check_mem(613,"000110101","001001010",0,'1'); -- (0, 0, 2, 1, 1, 2, 1, 2, 1)
sync_reset;
check_mem(614,"000110001","001001100",0,'1'); -- (0, 0, 2, 1, 1, 2, 2, 0, 1)
sync_reset;
check_mem(615,"000110010","001001100",1,'1'); -- (0, 0, 2, 1, 1, 2, 2, 1, 0)
sync_reset;
check_mem(616,"000110011","001001100",0,'1'); -- (0, 0, 2, 1, 1, 2, 2, 1, 1)
sync_reset;
check_mem(617,"000100001","001010000",6,'1'); -- (0, 0, 2, 1, 2, 0, 0, 0, 1)
sync_reset;
check_mem(618,"000100010","001010000",6,'1'); -- (0, 0, 2, 1, 2, 0, 0, 1, 0)
sync_reset;
check_mem(619,"000100011","001010000",6,'1'); -- (0, 0, 2, 1, 2, 0, 0, 1, 1)
sync_reset;
check_mem(620,"000100100","001010000",0,'1'); -- (0, 0, 2, 1, 2, 0, 1, 0, 0)
sync_reset;
check_mem(621,"000100101","001010000",0,'1'); -- (0, 0, 2, 1, 2, 0, 1, 0, 1)
sync_reset;
check_mem(622,"000100110","001010000",0,'1'); -- (0, 0, 2, 1, 2, 0, 1, 1, 0)
sync_reset;
check_mem(623,"000100110","001010001",0,'1'); -- (0, 0, 2, 1, 2, 0, 1, 1, 2)
sync_reset;
check_mem(624,"000100101","001010010",0,'1'); -- (0, 0, 2, 1, 2, 0, 1, 2, 1)
sync_reset;
check_mem(625,"000101000","001010000",0,'1'); -- (0, 0, 2, 1, 2, 1, 0, 0, 0)
sync_reset;
check_mem(626,"000101001","001010000",0,'1'); -- (0, 0, 2, 1, 2, 1, 0, 0, 1)
sync_reset;
check_mem(627,"000101010","001010000",0,'1'); -- (0, 0, 2, 1, 2, 1, 0, 1, 0)
sync_reset;
check_mem(628,"000101010","001010001",0,'1'); -- (0, 0, 2, 1, 2, 1, 0, 1, 2)
sync_reset;
check_mem(629,"000101001","001010010",0,'1'); -- (0, 0, 2, 1, 2, 1, 0, 2, 1)
sync_reset;
check_mem(630,"000101100","001010000",0,'1'); -- (0, 0, 2, 1, 2, 1, 1, 0, 0)
sync_reset;
check_mem(631,"000101100","001010001",0,'1'); -- (0, 0, 2, 1, 2, 1, 1, 0, 2)
sync_reset;
check_mem(632,"000101110","001010001",0,'1'); -- (0, 0, 2, 1, 2, 1, 1, 1, 2)
sync_reset;
check_mem(633,"000101100","001010010",0,'1'); -- (0, 0, 2, 1, 2, 1, 1, 2, 0)
sync_reset;
check_mem(634,"000101101","001010010",1,'1'); -- (0, 0, 2, 1, 2, 1, 1, 2, 1)
sync_reset;
check_mem(635,"000100011","001011000",6,'1'); -- (0, 0, 2, 1, 2, 2, 0, 1, 1)
sync_reset;
check_mem(636,"000100101","001011000",0,'1'); -- (0, 0, 2, 1, 2, 2, 1, 0, 1)
sync_reset;
check_mem(637,"000100110","001011000",0,'1'); -- (0, 0, 2, 1, 2, 2, 1, 1, 0)
sync_reset;
check_mem(638,"000000011","001100000",0,'1'); -- (0, 0, 2, 2, 0, 0, 0, 1, 1)
sync_reset;
check_mem(639,"000000101","001100000",0,'1'); -- (0, 0, 2, 2, 0, 0, 1, 0, 1)
sync_reset;
check_mem(640,"000000110","001100000",1,'1'); -- (0, 0, 2, 2, 0, 0, 1, 1, 0)
sync_reset;
check_mem(641,"000001001","001100000",0,'1'); -- (0, 0, 2, 2, 0, 1, 0, 0, 1)
sync_reset;
check_mem(642,"000001010","001100000",0,'1'); -- (0, 0, 2, 2, 0, 1, 0, 1, 0)
sync_reset;
check_mem(643,"000001011","001100000",6,'1'); -- (0, 0, 2, 2, 0, 1, 0, 1, 1)
sync_reset;
check_mem(644,"000001100","001100000",0,'1'); -- (0, 0, 2, 2, 0, 1, 1, 0, 0)
sync_reset;
check_mem(645,"000001101","001100000",7,'1'); -- (0, 0, 2, 2, 0, 1, 1, 0, 1)
sync_reset;
check_mem(646,"000001110","001100000",8,'1'); -- (0, 0, 2, 2, 0, 1, 1, 1, 0)
sync_reset;
check_mem(647,"000001110","001100001",0,'1'); -- (0, 0, 2, 2, 0, 1, 1, 1, 2)
sync_reset;
check_mem(648,"000001101","001100010",0,'1'); -- (0, 0, 2, 2, 0, 1, 1, 2, 1)
sync_reset;
check_mem(649,"000001011","001100100",0,'1'); -- (0, 0, 2, 2, 0, 1, 2, 1, 1)
sync_reset;
check_mem(650,"000010001","001100000",0,'1'); -- (0, 0, 2, 2, 1, 0, 0, 0, 1)
sync_reset;
check_mem(651,"000010010","001100000",0,'1'); -- (0, 0, 2, 2, 1, 0, 0, 1, 0)
sync_reset;
check_mem(652,"000010011","001100000",0,'1'); -- (0, 0, 2, 2, 1, 0, 0, 1, 1)
sync_reset;
check_mem(653,"000010100","001100000",7,'1'); -- (0, 0, 2, 2, 1, 0, 1, 0, 0)
sync_reset;
check_mem(654,"000010101","001100000",0,'1'); -- (0, 0, 2, 2, 1, 0, 1, 0, 1)
sync_reset;
check_mem(655,"000010110","001100000",0,'1'); -- (0, 0, 2, 2, 1, 0, 1, 1, 0)
sync_reset;
check_mem(656,"000010110","001100001",1,'1'); -- (0, 0, 2, 2, 1, 0, 1, 1, 2)
sync_reset;
check_mem(657,"000010101","001100010",0,'1'); -- (0, 0, 2, 2, 1, 0, 1, 2, 1)
sync_reset;
check_mem(658,"000010011","001100100",0,'1'); -- (0, 0, 2, 2, 1, 0, 2, 1, 1)
sync_reset;
check_mem(659,"000011000","001100000",0,'1'); -- (0, 0, 2, 2, 1, 1, 0, 0, 0)
sync_reset;
check_mem(660,"000011001","001100000",0,'1'); -- (0, 0, 2, 2, 1, 1, 0, 0, 1)
sync_reset;
check_mem(661,"000011010","001100000",1,'1'); -- (0, 0, 2, 2, 1, 1, 0, 1, 0)
sync_reset;
check_mem(662,"000011010","001100001",1,'1'); -- (0, 0, 2, 2, 1, 1, 0, 1, 2)
sync_reset;
check_mem(663,"000011001","001100010",0,'1'); -- (0, 0, 2, 2, 1, 1, 0, 2, 1)
sync_reset;
check_mem(664,"000011100","001100000",0,'1'); -- (0, 0, 2, 2, 1, 1, 1, 0, 0)
sync_reset;
check_mem(665,"000011100","001100001",0,'1'); -- (0, 0, 2, 2, 1, 1, 1, 0, 2)
sync_reset;
check_mem(666,"000011110","001100001",1,'1'); -- (0, 0, 2, 2, 1, 1, 1, 1, 2)
sync_reset;
check_mem(667,"000011100","001100010",0,'1'); -- (0, 0, 2, 2, 1, 1, 1, 2, 0)
sync_reset;
check_mem(668,"000011101","001100010",0,'1'); -- (0, 0, 2, 2, 1, 1, 1, 2, 1)
sync_reset;
check_mem(669,"000011001","001100100",0,'1'); -- (0, 0, 2, 2, 1, 1, 2, 0, 1)
sync_reset;
check_mem(670,"000011010","001100100",0,'1'); -- (0, 0, 2, 2, 1, 1, 2, 1, 0)
sync_reset;
check_mem(671,"000011011","001100100",0,'1'); -- (0, 0, 2, 2, 1, 1, 2, 1, 1)
sync_reset;
check_mem(672,"000010011","001101000",0,'1'); -- (0, 0, 2, 2, 1, 2, 0, 1, 1)
sync_reset;
check_mem(673,"000010101","001101000",0,'1'); -- (0, 0, 2, 2, 1, 2, 1, 0, 1)
sync_reset;
check_mem(674,"000010110","001101000",1,'1'); -- (0, 0, 2, 2, 1, 2, 1, 1, 0)
sync_reset;
check_mem(675,"000001011","001110000",6,'1'); -- (0, 0, 2, 2, 2, 1, 0, 1, 1)
sync_reset;
check_mem(676,"000001101","001110000",7,'1'); -- (0, 0, 2, 2, 2, 1, 1, 0, 1)
sync_reset;
check_mem(677,"000001110","001110000",8,'1'); -- (0, 0, 2, 2, 2, 1, 1, 1, 0)
sync_reset;
check_mem(678,"010000000","000000000",0,'1'); -- (0, 1, 0, 0, 0, 0, 0, 0, 0)
sync_reset;
check_mem(679,"010000000","000000001",2,'1'); -- (0, 1, 0, 0, 0, 0, 0, 0, 2)
sync_reset;
check_mem(680,"010000010","000000001",4,'1'); -- (0, 1, 0, 0, 0, 0, 0, 1, 2)
sync_reset;
check_mem(681,"010000000","000000010",0,'1'); -- (0, 1, 0, 0, 0, 0, 0, 2, 0)
sync_reset;
check_mem(682,"010000001","000000010",0,'1'); -- (0, 1, 0, 0, 0, 0, 0, 2, 1)
sync_reset;
check_mem(683,"010000100","000000001",2,'1'); -- (0, 1, 0, 0, 0, 0, 1, 0, 2)
sync_reset;
check_mem(684,"010000100","000000010",0,'1'); -- (0, 1, 0, 0, 0, 0, 1, 2, 0)
sync_reset;
check_mem(685,"010000100","000000011",0,'1'); -- (0, 1, 0, 0, 0, 0, 1, 2, 2)
sync_reset;
check_mem(686,"010000000","000000100",0,'1'); -- (0, 1, 0, 0, 0, 0, 2, 0, 0)
sync_reset;
check_mem(687,"010000001","000000100",0,'1'); -- (0, 1, 0, 0, 0, 0, 2, 0, 1)
sync_reset;
check_mem(688,"010000010","000000100",4,'1'); -- (0, 1, 0, 0, 0, 0, 2, 1, 0)
sync_reset;
check_mem(689,"010000010","000000101",0,'1'); -- (0, 1, 0, 0, 0, 0, 2, 1, 2)
sync_reset;
check_mem(690,"010000001","000000110",0,'1'); -- (0, 1, 0, 0, 0, 0, 2, 2, 1)
sync_reset;
check_mem(691,"010001000","000000001",6,'1'); -- (0, 1, 0, 0, 0, 1, 0, 0, 2)
sync_reset;
check_mem(692,"010001000","000000010",0,'1'); -- (0, 1, 0, 0, 0, 1, 0, 2, 0)
sync_reset;
check_mem(693,"010001000","000000011",6,'1'); -- (0, 1, 0, 0, 0, 1, 0, 2, 2)
sync_reset;
check_mem(694,"010001100","000000011",0,'1'); -- (0, 1, 0, 0, 0, 1, 1, 2, 2)
sync_reset;
check_mem(695,"010001000","000000100",0,'1'); -- (0, 1, 0, 0, 0, 1, 2, 0, 0)
sync_reset;
check_mem(696,"010001000","000000101",0,'1'); -- (0, 1, 0, 0, 0, 1, 2, 0, 2)
sync_reset;
check_mem(697,"010001010","000000101",4,'1'); -- (0, 1, 0, 0, 0, 1, 2, 1, 2)
sync_reset;
check_mem(698,"010001000","000000110",8,'1'); -- (0, 1, 0, 0, 0, 1, 2, 2, 0)
sync_reset;
check_mem(699,"010001001","000000110",0,'1'); -- (0, 1, 0, 0, 0, 1, 2, 2, 1)
sync_reset;
check_mem(700,"010000000","000001000",2,'1'); -- (0, 1, 0, 0, 0, 2, 0, 0, 0)
sync_reset;
check_mem(701,"010000001","000001000",4,'1'); -- (0, 1, 0, 0, 0, 2, 0, 0, 1)
sync_reset;
check_mem(702,"010000010","000001000",4,'1'); -- (0, 1, 0, 0, 0, 2, 0, 1, 0)
sync_reset;
check_mem(703,"010000010","000001001",2,'1'); -- (0, 1, 0, 0, 0, 2, 0, 1, 2)
sync_reset;
check_mem(704,"010000001","000001010",0,'1'); -- (0, 1, 0, 0, 0, 2, 0, 2, 1)
sync_reset;
check_mem(705,"010000100","000001000",4,'1'); -- (0, 1, 0, 0, 0, 2, 1, 0, 0)
sync_reset;
check_mem(706,"010000100","000001001",2,'1'); -- (0, 1, 0, 0, 0, 2, 1, 0, 2)
sync_reset;
check_mem(707,"010000110","000001001",2,'1'); -- (0, 1, 0, 0, 0, 2, 1, 1, 2)
sync_reset;
check_mem(708,"010000100","000001010",0,'1'); -- (0, 1, 0, 0, 0, 2, 1, 2, 0)
sync_reset;
check_mem(709,"010000101","000001010",0,'1'); -- (0, 1, 0, 0, 0, 2, 1, 2, 1)
sync_reset;
check_mem(710,"010000001","000001100",0,'1'); -- (0, 1, 0, 0, 0, 2, 2, 0, 1)
sync_reset;
check_mem(711,"010000010","000001100",0,'1'); -- (0, 1, 0, 0, 0, 2, 2, 1, 0)
sync_reset;
check_mem(712,"010000011","000001100",4,'1'); -- (0, 1, 0, 0, 0, 2, 2, 1, 1)
sync_reset;
check_mem(713,"010010000","000000001",7,'1'); -- (0, 1, 0, 0, 1, 0, 0, 0, 2)
sync_reset;
check_mem(714,"010010000","000000010",0,'1'); -- (0, 1, 0, 0, 1, 0, 0, 2, 0)
sync_reset;
check_mem(715,"010010000","000000011",6,'1'); -- (0, 1, 0, 0, 1, 0, 0, 2, 2)
sync_reset;
check_mem(716,"010010100","000000011",2,'1'); -- (0, 1, 0, 0, 1, 0, 1, 2, 2)
sync_reset;
check_mem(717,"010010000","000000100",7,'1'); -- (0, 1, 0, 0, 1, 0, 2, 0, 0)
sync_reset;
check_mem(718,"010010000","000000101",7,'1'); -- (0, 1, 0, 0, 1, 0, 2, 0, 2)
sync_reset;
check_mem(719,"010010000","000000110",8,'1'); -- (0, 1, 0, 0, 1, 0, 2, 2, 0)
sync_reset;
check_mem(720,"010010001","000000110",0,'1'); -- (0, 1, 0, 0, 1, 0, 2, 2, 1)
sync_reset;
check_mem(721,"010011000","000000011",6,'1'); -- (0, 1, 0, 0, 1, 1, 0, 2, 2)
sync_reset;
check_mem(722,"010011000","000000101",7,'1'); -- (0, 1, 0, 0, 1, 1, 2, 0, 2)
sync_reset;
check_mem(723,"010011000","000000110",3,'1'); -- (0, 1, 0, 0, 1, 1, 2, 2, 0)
sync_reset;
check_mem(724,"010010000","000001000",0,'1'); -- (0, 1, 0, 0, 1, 2, 0, 0, 0)
sync_reset;
check_mem(725,"010010000","000001001",2,'1'); -- (0, 1, 0, 0, 1, 2, 0, 0, 2)
sync_reset;
check_mem(726,"010010000","000001010",0,'1'); -- (0, 1, 0, 0, 1, 2, 0, 2, 0)
sync_reset;
check_mem(727,"010010001","000001010",0,'1'); -- (0, 1, 0, 0, 1, 2, 0, 2, 1)
sync_reset;
check_mem(728,"010010100","000001001",2,'1'); -- (0, 1, 0, 0, 1, 2, 1, 0, 2)
sync_reset;
check_mem(729,"010010100","000001010",2,'1'); -- (0, 1, 0, 0, 1, 2, 1, 2, 0)
sync_reset;
check_mem(730,"010010100","000001011",2,'1'); -- (0, 1, 0, 0, 1, 2, 1, 2, 2)
sync_reset;
check_mem(731,"010010000","000001100",0,'1'); -- (0, 1, 0, 0, 1, 2, 2, 0, 0)
sync_reset;
check_mem(732,"010010001","000001100",0,'1'); -- (0, 1, 0, 0, 1, 2, 2, 0, 1)
sync_reset;
check_mem(733,"010010001","000001110",0,'1'); -- (0, 1, 0, 0, 1, 2, 2, 2, 1)
sync_reset;
check_mem(734,"010000000","000010000",0,'1'); -- (0, 1, 0, 0, 2, 0, 0, 0, 0)
sync_reset;
check_mem(735,"010000001","000010000",0,'1'); -- (0, 1, 0, 0, 2, 0, 0, 0, 1)
sync_reset;
check_mem(736,"010000010","000010000",0,'1'); -- (0, 1, 0, 0, 2, 0, 0, 1, 0)
sync_reset;
check_mem(737,"010000010","000010001",0,'1'); -- (0, 1, 0, 0, 2, 0, 0, 1, 2)
sync_reset;
check_mem(738,"010000001","000010010",2,'1'); -- (0, 1, 0, 0, 2, 0, 0, 2, 1)
sync_reset;
check_mem(739,"010000100","000010000",0,'1'); -- (0, 1, 0, 0, 2, 0, 1, 0, 0)
sync_reset;
check_mem(740,"010000100","000010001",0,'1'); -- (0, 1, 0, 0, 2, 0, 1, 0, 2)
sync_reset;
check_mem(741,"010000110","000010001",0,'1'); -- (0, 1, 0, 0, 2, 0, 1, 1, 2)
sync_reset;
check_mem(742,"010000100","000010010",0,'1'); -- (0, 1, 0, 0, 2, 0, 1, 2, 0)
sync_reset;
check_mem(743,"010000101","000010010",0,'1'); -- (0, 1, 0, 0, 2, 0, 1, 2, 1)
sync_reset;
check_mem(744,"010000001","000010100",2,'1'); -- (0, 1, 0, 0, 2, 0, 2, 0, 1)
sync_reset;
check_mem(745,"010000010","000010100",0,'1'); -- (0, 1, 0, 0, 2, 0, 2, 1, 0)
sync_reset;
check_mem(746,"010000011","000010100",0,'1'); -- (0, 1, 0, 0, 2, 0, 2, 1, 1)
sync_reset;
check_mem(747,"010001000","000010000",0,'1'); -- (0, 1, 0, 0, 2, 1, 0, 0, 0)
sync_reset;
check_mem(748,"010001000","000010001",0,'1'); -- (0, 1, 0, 0, 2, 1, 0, 0, 2)
sync_reset;
check_mem(749,"010001010","000010001",0,'1'); -- (0, 1, 0, 0, 2, 1, 0, 1, 2)
sync_reset;
check_mem(750,"010001000","000010010",2,'1'); -- (0, 1, 0, 0, 2, 1, 0, 2, 0)
sync_reset;
check_mem(751,"010001001","000010010",2,'1'); -- (0, 1, 0, 0, 2, 1, 0, 2, 1)
sync_reset;
check_mem(752,"010001100","000010001",0,'1'); -- (0, 1, 0, 0, 2, 1, 1, 0, 2)
sync_reset;
check_mem(753,"010001100","000010010",0,'1'); -- (0, 1, 0, 0, 2, 1, 1, 2, 0)
sync_reset;
check_mem(754,"010001100","000010011",0,'1'); -- (0, 1, 0, 0, 2, 1, 1, 2, 2)
sync_reset;
check_mem(755,"010001000","000010100",2,'1'); -- (0, 1, 0, 0, 2, 1, 2, 0, 0)
sync_reset;
check_mem(756,"010001001","000010100",2,'1'); -- (0, 1, 0, 0, 2, 1, 2, 0, 1)
sync_reset;
check_mem(757,"010001010","000010100",0,'1'); -- (0, 1, 0, 0, 2, 1, 2, 1, 0)
sync_reset;
check_mem(758,"010001010","000010101",0,'1'); -- (0, 1, 0, 0, 2, 1, 2, 1, 2)
sync_reset;
check_mem(759,"010001001","000010110",2,'1'); -- (0, 1, 0, 0, 2, 1, 2, 2, 1)
sync_reset;
check_mem(760,"010000001","000011000",3,'1'); -- (0, 1, 0, 0, 2, 2, 0, 0, 1)
sync_reset;
check_mem(761,"010000010","000011000",0,'1'); -- (0, 1, 0, 0, 2, 2, 0, 1, 0)
sync_reset;
check_mem(762,"010000011","000011000",3,'1'); -- (0, 1, 0, 0, 2, 2, 0, 1, 1)
sync_reset;
check_mem(763,"010000100","000011000",3,'1'); -- (0, 1, 0, 0, 2, 2, 1, 0, 0)
sync_reset;
check_mem(764,"010000101","000011000",3,'1'); -- (0, 1, 0, 0, 2, 2, 1, 0, 1)
sync_reset;
check_mem(765,"010000110","000011000",3,'1'); -- (0, 1, 0, 0, 2, 2, 1, 1, 0)
sync_reset;
check_mem(766,"010000110","000011001",0,'1'); -- (0, 1, 0, 0, 2, 2, 1, 1, 2)
sync_reset;
check_mem(767,"010000101","000011010",3,'1'); -- (0, 1, 0, 0, 2, 2, 1, 2, 1)
sync_reset;
check_mem(768,"010000011","000011100",0,'1'); -- (0, 1, 0, 0, 2, 2, 2, 1, 1)
sync_reset;
check_mem(769,"010100000","000000001",2,'1'); -- (0, 1, 0, 1, 0, 0, 0, 0, 2)
sync_reset;
check_mem(770,"010100000","000000010",0,'1'); -- (0, 1, 0, 1, 0, 0, 0, 2, 0)
sync_reset;
check_mem(771,"010100000","000000011",6,'1'); -- (0, 1, 0, 1, 0, 0, 0, 2, 2)
sync_reset;
check_mem(772,"010100100","000000011",0,'1'); -- (0, 1, 0, 1, 0, 0, 1, 2, 2)
sync_reset;
check_mem(773,"010100000","000000100",8,'1'); -- (0, 1, 0, 1, 0, 0, 2, 0, 0)
sync_reset;
check_mem(774,"010100000","000000101",0,'1'); -- (0, 1, 0, 1, 0, 0, 2, 0, 2)
sync_reset;
check_mem(775,"010100010","000000101",4,'1'); -- (0, 1, 0, 1, 0, 0, 2, 1, 2)
sync_reset;
check_mem(776,"010100000","000000110",8,'1'); -- (0, 1, 0, 1, 0, 0, 2, 2, 0)
sync_reset;
check_mem(777,"010100001","000000110",0,'1'); -- (0, 1, 0, 1, 0, 0, 2, 2, 1)
sync_reset;
check_mem(778,"010101000","000000011",4,'1'); -- (0, 1, 0, 1, 0, 1, 0, 2, 2)
sync_reset;
check_mem(779,"010101000","000000101",4,'1'); -- (0, 1, 0, 1, 0, 1, 2, 0, 2)
sync_reset;
check_mem(780,"010101000","000000110",4,'1'); -- (0, 1, 0, 1, 0, 1, 2, 2, 0)
sync_reset;
check_mem(781,"010100000","000001000",0,'1'); -- (0, 1, 0, 1, 0, 2, 0, 0, 0)
sync_reset;
check_mem(782,"010100000","000001001",2,'1'); -- (0, 1, 0, 1, 0, 2, 0, 0, 2)
sync_reset;
check_mem(783,"010100010","000001001",2,'1'); -- (0, 1, 0, 1, 0, 2, 0, 1, 2)
sync_reset;
check_mem(784,"010100000","000001010",0,'1'); -- (0, 1, 0, 1, 0, 2, 0, 2, 0)
sync_reset;
check_mem(785,"010100001","000001010",0,'1'); -- (0, 1, 0, 1, 0, 2, 0, 2, 1)
sync_reset;
check_mem(786,"010100100","000001001",0,'1'); -- (0, 1, 0, 1, 0, 2, 1, 0, 2)
sync_reset;
check_mem(787,"010100100","000001010",0,'1'); -- (0, 1, 0, 1, 0, 2, 1, 2, 0)
sync_reset;
check_mem(788,"010100100","000001011",0,'1'); -- (0, 1, 0, 1, 0, 2, 1, 2, 2)
sync_reset;
check_mem(789,"010100000","000001100",2,'1'); -- (0, 1, 0, 1, 0, 2, 2, 0, 0)
sync_reset;
check_mem(790,"010100001","000001100",0,'1'); -- (0, 1, 0, 1, 0, 2, 2, 0, 1)
sync_reset;
check_mem(791,"010100010","000001100",4,'1'); -- (0, 1, 0, 1, 0, 2, 2, 1, 0)
sync_reset;
check_mem(792,"010100010","000001101",2,'1'); -- (0, 1, 0, 1, 0, 2, 2, 1, 2)
sync_reset;
check_mem(793,"010100001","000001110",0,'1'); -- (0, 1, 0, 1, 0, 2, 2, 2, 1)
sync_reset;
check_mem(794,"010110000","000000011",5,'1'); -- (0, 1, 0, 1, 1, 0, 0, 2, 2)
sync_reset;
check_mem(795,"010110000","000000101",7,'1'); -- (0, 1, 0, 1, 1, 0, 2, 0, 2)
sync_reset;
check_mem(796,"010110000","000000110",8,'1'); -- (0, 1, 0, 1, 1, 0, 2, 2, 0)
sync_reset;
check_mem(797,"010110000","000001001",2,'1'); -- (0, 1, 0, 1, 1, 2, 0, 0, 2)
sync_reset;
check_mem(798,"010110000","000001010",8,'1'); -- (0, 1, 0, 1, 1, 2, 0, 2, 0)
sync_reset;
check_mem(799,"010110000","000001011",0,'1'); -- (0, 1, 0, 1, 1, 2, 0, 2, 2)
sync_reset;
check_mem(800,"010110100","000001011",2,'1'); -- (0, 1, 0, 1, 1, 2, 1, 2, 2)
sync_reset;
check_mem(801,"010110000","000001100",7,'1'); -- (0, 1, 0, 1, 1, 2, 2, 0, 0)
sync_reset;
check_mem(802,"010110000","000001101",7,'1'); -- (0, 1, 0, 1, 1, 2, 2, 0, 2)
sync_reset;
check_mem(803,"010110000","000001110",8,'1'); -- (0, 1, 0, 1, 1, 2, 2, 2, 0)
sync_reset;
check_mem(804,"010110001","000001110",0,'1'); -- (0, 1, 0, 1, 1, 2, 2, 2, 1)
sync_reset;
check_mem(805,"010100000","000010000",0,'1'); -- (0, 1, 0, 1, 2, 0, 0, 0, 0)
sync_reset;
check_mem(806,"010100000","000010001",0,'1'); -- (0, 1, 0, 1, 2, 0, 0, 0, 2)
sync_reset;
check_mem(807,"010100010","000010001",0,'1'); -- (0, 1, 0, 1, 2, 0, 0, 1, 2)
sync_reset;
check_mem(808,"010100000","000010010",0,'1'); -- (0, 1, 0, 1, 2, 0, 0, 2, 0)
sync_reset;
check_mem(809,"010100001","000010010",0,'1'); -- (0, 1, 0, 1, 2, 0, 0, 2, 1)
sync_reset;
check_mem(810,"010100100","000010001",0,'1'); -- (0, 1, 0, 1, 2, 0, 1, 0, 2)
sync_reset;
check_mem(811,"010100100","000010010",0,'1'); -- (0, 1, 0, 1, 2, 0, 1, 2, 0)
sync_reset;
check_mem(812,"010100100","000010011",0,'1'); -- (0, 1, 0, 1, 2, 0, 1, 2, 2)
sync_reset;
check_mem(813,"010100000","000010100",2,'1'); -- (0, 1, 0, 1, 2, 0, 2, 0, 0)
sync_reset;
check_mem(814,"010100001","000010100",2,'1'); -- (0, 1, 0, 1, 2, 0, 2, 0, 1)
sync_reset;
check_mem(815,"010100010","000010100",0,'1'); -- (0, 1, 0, 1, 2, 0, 2, 1, 0)
sync_reset;
check_mem(816,"010100010","000010101",0,'1'); -- (0, 1, 0, 1, 2, 0, 2, 1, 2)
sync_reset;
check_mem(817,"010100001","000010110",2,'1'); -- (0, 1, 0, 1, 2, 0, 2, 2, 1)
sync_reset;
check_mem(818,"010101000","000010001",0,'1'); -- (0, 1, 0, 1, 2, 1, 0, 0, 2)
sync_reset;
check_mem(819,"010101000","000010010",6,'1'); -- (0, 1, 0, 1, 2, 1, 0, 2, 0)
sync_reset;
check_mem(820,"010101000","000010011",0,'1'); -- (0, 1, 0, 1, 2, 1, 0, 2, 2)
sync_reset;
check_mem(821,"010101100","000010011",0,'1'); -- (0, 1, 0, 1, 2, 1, 1, 2, 2)
sync_reset;
check_mem(822,"010101000","000010100",0,'1'); -- (0, 1, 0, 1, 2, 1, 2, 0, 0)
sync_reset;
check_mem(823,"010101000","000010101",0,'1'); -- (0, 1, 0, 1, 2, 1, 2, 0, 2)
sync_reset;
check_mem(824,"010101010","000010101",0,'1'); -- (0, 1, 0, 1, 2, 1, 2, 1, 2)
sync_reset;
check_mem(825,"010101000","000010110",0,'1'); -- (0, 1, 0, 1, 2, 1, 2, 2, 0)
sync_reset;
check_mem(826,"010101001","000010110",2,'1'); -- (0, 1, 0, 1, 2, 1, 2, 2, 1)
sync_reset;
check_mem(827,"010100000","000011000",0,'1'); -- (0, 1, 0, 1, 2, 2, 0, 0, 0)
sync_reset;
check_mem(828,"010100001","000011000",0,'1'); -- (0, 1, 0, 1, 2, 2, 0, 0, 1)
sync_reset;
check_mem(829,"010100010","000011000",2,'1'); -- (0, 1, 0, 1, 2, 2, 0, 1, 0)
sync_reset;
check_mem(830,"010100010","000011001",0,'1'); -- (0, 1, 0, 1, 2, 2, 0, 1, 2)
sync_reset;
check_mem(831,"010100001","000011010",0,'1'); -- (0, 1, 0, 1, 2, 2, 0, 2, 1)
sync_reset;
check_mem(832,"010100100","000011000",0,'1'); -- (0, 1, 0, 1, 2, 2, 1, 0, 0)
sync_reset;
check_mem(833,"010100100","000011001",0,'1'); -- (0, 1, 0, 1, 2, 2, 1, 0, 2)
sync_reset;
check_mem(834,"010100110","000011001",0,'1'); -- (0, 1, 0, 1, 2, 2, 1, 1, 2)
sync_reset;
check_mem(835,"010100100","000011010",0,'1'); -- (0, 1, 0, 1, 2, 2, 1, 2, 0)
sync_reset;
check_mem(836,"010100101","000011010",0,'1'); -- (0, 1, 0, 1, 2, 2, 1, 2, 1)
sync_reset;
check_mem(837,"010100001","000011100",2,'1'); -- (0, 1, 0, 1, 2, 2, 2, 0, 1)
sync_reset;
check_mem(838,"010100010","000011100",2,'1'); -- (0, 1, 0, 1, 2, 2, 2, 1, 0)
sync_reset;
check_mem(839,"010100011","000011100",2,'1'); -- (0, 1, 0, 1, 2, 2, 2, 1, 1)
sync_reset;
check_mem(840,"010000000","000100000",0,'1'); -- (0, 1, 0, 2, 0, 0, 0, 0, 0)
sync_reset;
check_mem(841,"010000001","000100000",4,'1'); -- (0, 1, 0, 2, 0, 0, 0, 0, 1)
sync_reset;
check_mem(842,"010000010","000100000",4,'1'); -- (0, 1, 0, 2, 0, 0, 0, 1, 0)
sync_reset;
check_mem(843,"010000010","000100001",0,'1'); -- (0, 1, 0, 2, 0, 0, 0, 1, 2)
sync_reset;
check_mem(844,"010000001","000100010",0,'1'); -- (0, 1, 0, 2, 0, 0, 0, 2, 1)
sync_reset;
check_mem(845,"010000100","000100000",4,'1'); -- (0, 1, 0, 2, 0, 0, 1, 0, 0)
sync_reset;
check_mem(846,"010000100","000100001",2,'1'); -- (0, 1, 0, 2, 0, 0, 1, 0, 2)
sync_reset;
check_mem(847,"010000110","000100001",4,'1'); -- (0, 1, 0, 2, 0, 0, 1, 1, 2)
sync_reset;
check_mem(848,"010000100","000100010",2,'1'); -- (0, 1, 0, 2, 0, 0, 1, 2, 0)
sync_reset;
check_mem(849,"010000101","000100010",2,'1'); -- (0, 1, 0, 2, 0, 0, 1, 2, 1)
sync_reset;
check_mem(850,"010000001","000100100",0,'1'); -- (0, 1, 0, 2, 0, 0, 2, 0, 1)
sync_reset;
check_mem(851,"010000010","000100100",0,'1'); -- (0, 1, 0, 2, 0, 0, 2, 1, 0)
sync_reset;
check_mem(852,"010000011","000100100",0,'1'); -- (0, 1, 0, 2, 0, 0, 2, 1, 1)
sync_reset;
check_mem(853,"010001000","000100000",2,'1'); -- (0, 1, 0, 2, 0, 1, 0, 0, 0)
sync_reset;
check_mem(854,"010001000","000100001",0,'1'); -- (0, 1, 0, 2, 0, 1, 0, 0, 2)
sync_reset;
check_mem(855,"010001010","000100001",4,'1'); -- (0, 1, 0, 2, 0, 1, 0, 1, 2)
sync_reset;
check_mem(856,"010001000","000100010",2,'1'); -- (0, 1, 0, 2, 0, 1, 0, 2, 0)
sync_reset;
check_mem(857,"010001001","000100010",2,'1'); -- (0, 1, 0, 2, 0, 1, 0, 2, 1)
sync_reset;
check_mem(858,"010001100","000100001",2,'1'); -- (0, 1, 0, 2, 0, 1, 1, 0, 2)
sync_reset;
check_mem(859,"010001100","000100010",2,'1'); -- (0, 1, 0, 2, 0, 1, 1, 2, 0)
sync_reset;
check_mem(860,"010001100","000100011",2,'1'); -- (0, 1, 0, 2, 0, 1, 1, 2, 2)
sync_reset;
check_mem(861,"010001000","000100100",0,'1'); -- (0, 1, 0, 2, 0, 1, 2, 0, 0)
sync_reset;
check_mem(862,"010001001","000100100",0,'1'); -- (0, 1, 0, 2, 0, 1, 2, 0, 1)
sync_reset;
check_mem(863,"010001010","000100100",0,'1'); -- (0, 1, 0, 2, 0, 1, 2, 1, 0)
sync_reset;
check_mem(864,"010001010","000100101",0,'1'); -- (0, 1, 0, 2, 0, 1, 2, 1, 2)
sync_reset;
check_mem(865,"010001001","000100110",0,'1'); -- (0, 1, 0, 2, 0, 1, 2, 2, 1)
sync_reset;
check_mem(866,"010000001","000101000",4,'1'); -- (0, 1, 0, 2, 0, 2, 0, 0, 1)
sync_reset;
check_mem(867,"010000010","000101000",4,'1'); -- (0, 1, 0, 2, 0, 2, 0, 1, 0)
sync_reset;
check_mem(868,"010000011","000101000",4,'1'); -- (0, 1, 0, 2, 0, 2, 0, 1, 1)
sync_reset;
check_mem(869,"010000100","000101000",4,'1'); -- (0, 1, 0, 2, 0, 2, 1, 0, 0)
sync_reset;
check_mem(870,"010000101","000101000",4,'1'); -- (0, 1, 0, 2, 0, 2, 1, 0, 1)
sync_reset;
check_mem(871,"010000110","000101000",4,'1'); -- (0, 1, 0, 2, 0, 2, 1, 1, 0)
sync_reset;
check_mem(872,"010000110","000101001",4,'1'); -- (0, 1, 0, 2, 0, 2, 1, 1, 2)
sync_reset;
check_mem(873,"010000101","000101010",4,'1'); -- (0, 1, 0, 2, 0, 2, 1, 2, 1)
sync_reset;
check_mem(874,"010000011","000101100",4,'1'); -- (0, 1, 0, 2, 0, 2, 2, 1, 1)
sync_reset;
check_mem(875,"010010000","000100000",0,'1'); -- (0, 1, 0, 2, 1, 0, 0, 0, 0)
sync_reset;
check_mem(876,"010010000","000100001",0,'1'); -- (0, 1, 0, 2, 1, 0, 0, 0, 2)
sync_reset;
check_mem(877,"010010000","000100010",0,'1'); -- (0, 1, 0, 2, 1, 0, 0, 2, 0)
sync_reset;
check_mem(878,"010010001","000100010",0,'1'); -- (0, 1, 0, 2, 1, 0, 0, 2, 1)
sync_reset;
check_mem(879,"010010100","000100001",0,'1'); -- (0, 1, 0, 2, 1, 0, 1, 0, 2)
sync_reset;
check_mem(880,"010010100","000100010",2,'1'); -- (0, 1, 0, 2, 1, 0, 1, 2, 0)
sync_reset;
check_mem(881,"010010100","000100011",2,'1'); -- (0, 1, 0, 2, 1, 0, 1, 2, 2)
sync_reset;
check_mem(882,"010010000","000100100",0,'1'); -- (0, 1, 0, 2, 1, 0, 2, 0, 0)
sync_reset;
check_mem(883,"010010001","000100100",0,'1'); -- (0, 1, 0, 2, 1, 0, 2, 0, 1)
sync_reset;
check_mem(884,"010010001","000100110",0,'1'); -- (0, 1, 0, 2, 1, 0, 2, 2, 1)
sync_reset;
check_mem(885,"010011000","000100001",7,'1'); -- (0, 1, 0, 2, 1, 1, 0, 0, 2)
sync_reset;
check_mem(886,"010011000","000100010",6,'1'); -- (0, 1, 0, 2, 1, 1, 0, 2, 0)
sync_reset;
check_mem(887,"010011000","000100011",6,'1'); -- (0, 1, 0, 2, 1, 1, 0, 2, 2)
sync_reset;
check_mem(888,"010011100","000100011",2,'1'); -- (0, 1, 0, 2, 1, 1, 1, 2, 2)
sync_reset;
check_mem(889,"010011000","000100100",0,'1'); -- (0, 1, 0, 2, 1, 1, 2, 0, 0)
sync_reset;
check_mem(890,"010011000","000100101",7,'1'); -- (0, 1, 0, 2, 1, 1, 2, 0, 2)
sync_reset;
check_mem(891,"010011000","000100110",0,'1'); -- (0, 1, 0, 2, 1, 1, 2, 2, 0)
sync_reset;
check_mem(892,"010011001","000100110",0,'1'); -- (0, 1, 0, 2, 1, 1, 2, 2, 1)
sync_reset;
check_mem(893,"010010000","000101000",0,'1'); -- (0, 1, 0, 2, 1, 2, 0, 0, 0)
sync_reset;
check_mem(894,"010010001","000101000",0,'1'); -- (0, 1, 0, 2, 1, 2, 0, 0, 1)
sync_reset;
check_mem(895,"010010001","000101010",0,'1'); -- (0, 1, 0, 2, 1, 2, 0, 2, 1)
sync_reset;
check_mem(896,"010010100","000101000",0,'1'); -- (0, 1, 0, 2, 1, 2, 1, 0, 0)
sync_reset;
check_mem(897,"010010100","000101001",2,'1'); -- (0, 1, 0, 2, 1, 2, 1, 0, 2)
sync_reset;
check_mem(898,"010010100","000101010",0,'1'); -- (0, 1, 0, 2, 1, 2, 1, 2, 0)
sync_reset;
check_mem(899,"010010101","000101010",0,'1'); -- (0, 1, 0, 2, 1, 2, 1, 2, 1)
sync_reset;
check_mem(900,"010010001","000101100",0,'1'); -- (0, 1, 0, 2, 1, 2, 2, 0, 1)
sync_reset;
check_mem(901,"010000001","000110000",5,'1'); -- (0, 1, 0, 2, 2, 0, 0, 0, 1)
sync_reset;
check_mem(902,"010000010","000110000",0,'1'); -- (0, 1, 0, 2, 2, 0, 0, 1, 0)
sync_reset;
check_mem(903,"010000011","000110000",5,'1'); -- (0, 1, 0, 2, 2, 0, 0, 1, 1)
sync_reset;
check_mem(904,"010000100","000110000",5,'1'); -- (0, 1, 0, 2, 2, 0, 1, 0, 0)
sync_reset;
check_mem(905,"010000101","000110000",5,'1'); -- (0, 1, 0, 2, 2, 0, 1, 0, 1)
sync_reset;
check_mem(906,"010000110","000110000",5,'1'); -- (0, 1, 0, 2, 2, 0, 1, 1, 0)
sync_reset;
check_mem(907,"010000110","000110001",0,'1'); -- (0, 1, 0, 2, 2, 0, 1, 1, 2)
sync_reset;
check_mem(908,"010000101","000110010",5,'1'); -- (0, 1, 0, 2, 2, 0, 1, 2, 1)
sync_reset;
check_mem(909,"010000011","000110100",0,'1'); -- (0, 1, 0, 2, 2, 0, 2, 1, 1)
sync_reset;
check_mem(910,"010001000","000110000",2,'1'); -- (0, 1, 0, 2, 2, 1, 0, 0, 0)
sync_reset;
check_mem(911,"010001001","000110000",2,'1'); -- (0, 1, 0, 2, 2, 1, 0, 0, 1)
sync_reset;
check_mem(912,"010001010","000110000",0,'1'); -- (0, 1, 0, 2, 2, 1, 0, 1, 0)
sync_reset;
check_mem(913,"010001010","000110001",0,'1'); -- (0, 1, 0, 2, 2, 1, 0, 1, 2)
sync_reset;
check_mem(914,"010001001","000110010",2,'1'); -- (0, 1, 0, 2, 2, 1, 0, 2, 1)
sync_reset;
check_mem(915,"010001100","000110000",2,'1'); -- (0, 1, 0, 2, 2, 1, 1, 0, 0)
sync_reset;
check_mem(916,"010001100","000110001",0,'1'); -- (0, 1, 0, 2, 2, 1, 1, 0, 2)
sync_reset;
check_mem(917,"010001110","000110001",0,'1'); -- (0, 1, 0, 2, 2, 1, 1, 1, 2)
sync_reset;
check_mem(918,"010001100","000110010",2,'1'); -- (0, 1, 0, 2, 2, 1, 1, 2, 0)
sync_reset;
check_mem(919,"010001101","000110010",2,'1'); -- (0, 1, 0, 2, 2, 1, 1, 2, 1)
sync_reset;
check_mem(920,"010001001","000110100",2,'1'); -- (0, 1, 0, 2, 2, 1, 2, 0, 1)
sync_reset;
check_mem(921,"010001010","000110100",0,'1'); -- (0, 1, 0, 2, 2, 1, 2, 1, 0)
sync_reset;
check_mem(922,"010001011","000110100",0,'1'); -- (0, 1, 0, 2, 2, 1, 2, 1, 1)
sync_reset;
check_mem(923,"011000000","000000001",0,'1'); -- (0, 1, 1, 0, 0, 0, 0, 0, 2)
sync_reset;
check_mem(924,"011000000","000000010",0,'1'); -- (0, 1, 1, 0, 0, 0, 0, 2, 0)
sync_reset;
check_mem(925,"011000000","000000011",0,'1'); -- (0, 1, 1, 0, 0, 0, 0, 2, 2)
sync_reset;
check_mem(926,"011000100","000000011",0,'1'); -- (0, 1, 1, 0, 0, 0, 1, 2, 2)
sync_reset;
check_mem(927,"011000000","000000100",0,'1'); -- (0, 1, 1, 0, 0, 0, 2, 0, 0)
sync_reset;
check_mem(928,"011000000","000000101",0,'1'); -- (0, 1, 1, 0, 0, 0, 2, 0, 2)
sync_reset;
check_mem(929,"011000010","000000101",0,'1'); -- (0, 1, 1, 0, 0, 0, 2, 1, 2)
sync_reset;
check_mem(930,"011000000","000000110",0,'1'); -- (0, 1, 1, 0, 0, 0, 2, 2, 0)
sync_reset;
check_mem(931,"011000001","000000110",0,'1'); -- (0, 1, 1, 0, 0, 0, 2, 2, 1)
sync_reset;
check_mem(932,"011001000","000000011",0,'1'); -- (0, 1, 1, 0, 0, 1, 0, 2, 2)
sync_reset;
check_mem(933,"011001000","000000101",0,'1'); -- (0, 1, 1, 0, 0, 1, 2, 0, 2)
sync_reset;
check_mem(934,"011001000","000000110",8,'1'); -- (0, 1, 1, 0, 0, 1, 2, 2, 0)
sync_reset;
check_mem(935,"011000000","000001000",0,'1'); -- (0, 1, 1, 0, 0, 2, 0, 0, 0)
sync_reset;
check_mem(936,"011000000","000001001",0,'1'); -- (0, 1, 1, 0, 0, 2, 0, 0, 2)
sync_reset;
check_mem(937,"011000010","000001001",0,'1'); -- (0, 1, 1, 0, 0, 2, 0, 1, 2)
sync_reset;
check_mem(938,"011000000","000001010",0,'1'); -- (0, 1, 1, 0, 0, 2, 0, 2, 0)
sync_reset;
check_mem(939,"011000001","000001010",0,'1'); -- (0, 1, 1, 0, 0, 2, 0, 2, 1)
sync_reset;
check_mem(940,"011000100","000001001",0,'1'); -- (0, 1, 1, 0, 0, 2, 1, 0, 2)
sync_reset;
check_mem(941,"011000100","000001010",0,'1'); -- (0, 1, 1, 0, 0, 2, 1, 2, 0)
sync_reset;
check_mem(942,"011000100","000001011",0,'1'); -- (0, 1, 1, 0, 0, 2, 1, 2, 2)
sync_reset;
check_mem(943,"011000000","000001100",0,'1'); -- (0, 1, 1, 0, 0, 2, 2, 0, 0)
sync_reset;
check_mem(944,"011000001","000001100",0,'1'); -- (0, 1, 1, 0, 0, 2, 2, 0, 1)
sync_reset;
check_mem(945,"011000010","000001100",0,'1'); -- (0, 1, 1, 0, 0, 2, 2, 1, 0)
sync_reset;
check_mem(946,"011000010","000001101",0,'1'); -- (0, 1, 1, 0, 0, 2, 2, 1, 2)
sync_reset;
check_mem(947,"011000001","000001110",0,'1'); -- (0, 1, 1, 0, 0, 2, 2, 2, 1)
sync_reset;
check_mem(948,"011010000","000000011",6,'1'); -- (0, 1, 1, 0, 1, 0, 0, 2, 2)
sync_reset;
check_mem(949,"011010000","000000101",7,'1'); -- (0, 1, 1, 0, 1, 0, 2, 0, 2)
sync_reset;
check_mem(950,"011010000","000000110",0,'1'); -- (0, 1, 1, 0, 1, 0, 2, 2, 0)
sync_reset;
check_mem(951,"011010000","000001001",0,'1'); -- (0, 1, 1, 0, 1, 2, 0, 0, 2)
sync_reset;
check_mem(952,"011010000","000001010",0,'1'); -- (0, 1, 1, 0, 1, 2, 0, 2, 0)
sync_reset;
check_mem(953,"011010000","000001011",0,'1'); -- (0, 1, 1, 0, 1, 2, 0, 2, 2)
sync_reset;
check_mem(954,"011010000","000001100",0,'1'); -- (0, 1, 1, 0, 1, 2, 2, 0, 0)
sync_reset;
check_mem(955,"011010000","000001101",0,'1'); -- (0, 1, 1, 0, 1, 2, 2, 0, 2)
sync_reset;
check_mem(956,"011010000","000001110",0,'1'); -- (0, 1, 1, 0, 1, 2, 2, 2, 0)
sync_reset;
check_mem(957,"011010001","000001110",0,'1'); -- (0, 1, 1, 0, 1, 2, 2, 2, 1)
sync_reset;
check_mem(958,"011000000","000010000",0,'1'); -- (0, 1, 1, 0, 2, 0, 0, 0, 0)
sync_reset;
check_mem(959,"011000000","000010001",0,'1'); -- (0, 1, 1, 0, 2, 0, 0, 0, 2)
sync_reset;
check_mem(960,"011000010","000010001",0,'1'); -- (0, 1, 1, 0, 2, 0, 0, 1, 2)
sync_reset;
check_mem(961,"011000000","000010010",0,'1'); -- (0, 1, 1, 0, 2, 0, 0, 2, 0)
sync_reset;
check_mem(962,"011000001","000010010",0,'1'); -- (0, 1, 1, 0, 2, 0, 0, 2, 1)
sync_reset;
check_mem(963,"011000100","000010001",0,'1'); -- (0, 1, 1, 0, 2, 0, 1, 0, 2)
sync_reset;
check_mem(964,"011000100","000010010",0,'1'); -- (0, 1, 1, 0, 2, 0, 1, 2, 0)
sync_reset;
check_mem(965,"011000100","000010011",0,'1'); -- (0, 1, 1, 0, 2, 0, 1, 2, 2)
sync_reset;
check_mem(966,"011000000","000010100",0,'1'); -- (0, 1, 1, 0, 2, 0, 2, 0, 0)
sync_reset;
check_mem(967,"011000001","000010100",0,'1'); -- (0, 1, 1, 0, 2, 0, 2, 0, 1)
sync_reset;
check_mem(968,"011000010","000010100",0,'1'); -- (0, 1, 1, 0, 2, 0, 2, 1, 0)
sync_reset;
check_mem(969,"011000010","000010101",0,'1'); -- (0, 1, 1, 0, 2, 0, 2, 1, 2)
sync_reset;
check_mem(970,"011000001","000010110",0,'1'); -- (0, 1, 1, 0, 2, 0, 2, 2, 1)
sync_reset;
check_mem(971,"011001000","000010001",0,'1'); -- (0, 1, 1, 0, 2, 1, 0, 0, 2)
sync_reset;
check_mem(972,"011001000","000010010",0,'1'); -- (0, 1, 1, 0, 2, 1, 0, 2, 0)
sync_reset;
check_mem(973,"011001000","000010011",0,'1'); -- (0, 1, 1, 0, 2, 1, 0, 2, 2)
sync_reset;
check_mem(974,"011001100","000010011",0,'1'); -- (0, 1, 1, 0, 2, 1, 1, 2, 2)
sync_reset;
check_mem(975,"011001000","000010100",0,'1'); -- (0, 1, 1, 0, 2, 1, 2, 0, 0)
sync_reset;
check_mem(976,"011001000","000010101",0,'1'); -- (0, 1, 1, 0, 2, 1, 2, 0, 2)
sync_reset;
check_mem(977,"011001010","000010101",0,'1'); -- (0, 1, 1, 0, 2, 1, 2, 1, 2)
sync_reset;
check_mem(978,"011001000","000010110",0,'1'); -- (0, 1, 1, 0, 2, 1, 2, 2, 0)
sync_reset;
check_mem(979,"011000000","000011000",0,'1'); -- (0, 1, 1, 0, 2, 2, 0, 0, 0)
sync_reset;
check_mem(980,"011000001","000011000",3,'1'); -- (0, 1, 1, 0, 2, 2, 0, 0, 1)
sync_reset;
check_mem(981,"011000010","000011000",0,'1'); -- (0, 1, 1, 0, 2, 2, 0, 1, 0)
sync_reset;
check_mem(982,"011000010","000011001",0,'1'); -- (0, 1, 1, 0, 2, 2, 0, 1, 2)
sync_reset;
check_mem(983,"011000001","000011010",0,'1'); -- (0, 1, 1, 0, 2, 2, 0, 2, 1)
sync_reset;
check_mem(984,"011000100","000011000",0,'1'); -- (0, 1, 1, 0, 2, 2, 1, 0, 0)
sync_reset;
check_mem(985,"011000100","000011001",0,'1'); -- (0, 1, 1, 0, 2, 2, 1, 0, 2)
sync_reset;
check_mem(986,"011000110","000011001",0,'1'); -- (0, 1, 1, 0, 2, 2, 1, 1, 2)
sync_reset;
check_mem(987,"011000100","000011010",0,'1'); -- (0, 1, 1, 0, 2, 2, 1, 2, 0)
sync_reset;
check_mem(988,"011000101","000011010",3,'1'); -- (0, 1, 1, 0, 2, 2, 1, 2, 1)
sync_reset;
check_mem(989,"011000001","000011100",0,'1'); -- (0, 1, 1, 0, 2, 2, 2, 0, 1)
sync_reset;
check_mem(990,"011000010","000011100",0,'1'); -- (0, 1, 1, 0, 2, 2, 2, 1, 0)
sync_reset;
check_mem(991,"011000011","000011100",3,'1'); -- (0, 1, 1, 0, 2, 2, 2, 1, 1)
sync_reset;
check_mem(992,"011100000","000000011",0,'1'); -- (0, 1, 1, 1, 0, 0, 0, 2, 2)
sync_reset;
check_mem(993,"011100000","000000101",0,'1'); -- (0, 1, 1, 1, 0, 0, 2, 0, 2)
sync_reset;
check_mem(994,"011100000","000000110",8,'1'); -- (0, 1, 1, 1, 0, 0, 2, 2, 0)
sync_reset;
check_mem(995,"011100000","000001001",0,'1'); -- (0, 1, 1, 1, 0, 2, 0, 0, 2)
sync_reset;
check_mem(996,"011100000","000001010",0,'1'); -- (0, 1, 1, 1, 0, 2, 0, 2, 0)
sync_reset;
check_mem(997,"011100000","000001011",0,'1'); -- (0, 1, 1, 1, 0, 2, 0, 2, 2)
sync_reset;
check_mem(998,"011100100","000001011",0,'1'); -- (0, 1, 1, 1, 0, 2, 1, 2, 2)
sync_reset;
check_mem(999,"011100000","000001100",0,'1'); -- (0, 1, 1, 1, 0, 2, 2, 0, 0)
sync_reset;
check_mem(1000,"011100000","000001101",0,'1'); -- (0, 1, 1, 1, 0, 2, 2, 0, 2)
sync_reset;
check_mem(1001,"011100010","000001101",0,'1'); -- (0, 1, 1, 1, 0, 2, 2, 1, 2)
sync_reset;
check_mem(1002,"011100000","000001110",0,'1'); -- (0, 1, 1, 1, 0, 2, 2, 2, 0)
sync_reset;
check_mem(1003,"011100001","000001110",0,'1'); -- (0, 1, 1, 1, 0, 2, 2, 2, 1)
sync_reset;
check_mem(1004,"011110000","000001011",6,'1'); -- (0, 1, 1, 1, 1, 2, 0, 2, 2)
sync_reset;
check_mem(1005,"011110000","000001101",7,'1'); -- (0, 1, 1, 1, 1, 2, 2, 0, 2)
sync_reset;
check_mem(1006,"011110000","000001110",8,'1'); -- (0, 1, 1, 1, 1, 2, 2, 2, 0)
sync_reset;
check_mem(1007,"011100000","000010001",0,'1'); -- (0, 1, 1, 1, 2, 0, 0, 0, 2)
sync_reset;
check_mem(1008,"011100000","000010010",0,'1'); -- (0, 1, 1, 1, 2, 0, 0, 2, 0)
sync_reset;
check_mem(1009,"011100000","000010011",0,'1'); -- (0, 1, 1, 1, 2, 0, 0, 2, 2)
sync_reset;
check_mem(1010,"011100100","000010011",0,'1'); -- (0, 1, 1, 1, 2, 0, 1, 2, 2)
sync_reset;
check_mem(1011,"011100000","000010100",0,'1'); -- (0, 1, 1, 1, 2, 0, 2, 0, 0)
sync_reset;
check_mem(1012,"011100000","000010101",0,'1'); -- (0, 1, 1, 1, 2, 0, 2, 0, 2)
sync_reset;
check_mem(1013,"011100010","000010101",0,'1'); -- (0, 1, 1, 1, 2, 0, 2, 1, 2)
sync_reset;
check_mem(1014,"011100000","000010110",0,'1'); -- (0, 1, 1, 1, 2, 0, 2, 2, 0)
sync_reset;
check_mem(1015,"011100001","000010110",0,'1'); -- (0, 1, 1, 1, 2, 0, 2, 2, 1)
sync_reset;
check_mem(1016,"011101000","000010011",0,'1'); -- (0, 1, 1, 1, 2, 1, 0, 2, 2)
sync_reset;
check_mem(1017,"011101000","000010101",0,'1'); -- (0, 1, 1, 1, 2, 1, 2, 0, 2)
sync_reset;
check_mem(1018,"011101000","000010110",8,'1'); -- (0, 1, 1, 1, 2, 1, 2, 2, 0)
sync_reset;
check_mem(1019,"011100000","000011000",0,'1'); -- (0, 1, 1, 1, 2, 2, 0, 0, 0)
sync_reset;
check_mem(1020,"011100000","000011001",0,'1'); -- (0, 1, 1, 1, 2, 2, 0, 0, 2)
sync_reset;
check_mem(1021,"011100010","000011001",0,'1'); -- (0, 1, 1, 1, 2, 2, 0, 1, 2)
sync_reset;
check_mem(1022,"011100000","000011010",0,'1'); -- (0, 1, 1, 1, 2, 2, 0, 2, 0)
sync_reset;
check_mem(1023,"011100001","000011010",0,'1'); -- (0, 1, 1, 1, 2, 2, 0, 2, 1)
sync_reset;
check_mem(1024,"011100100","000011001",0,'1'); -- (0, 1, 1, 1, 2, 2, 1, 0, 2)
sync_reset;
check_mem(1025,"011100100","000011010",0,'1'); -- (0, 1, 1, 1, 2, 2, 1, 2, 0)
sync_reset;
check_mem(1026,"011100100","000011011",0,'1'); -- (0, 1, 1, 1, 2, 2, 1, 2, 2)
sync_reset;
check_mem(1027,"011100000","000011100",0,'1'); -- (0, 1, 1, 1, 2, 2, 2, 0, 0)
sync_reset;
check_mem(1028,"011100001","000011100",0,'1'); -- (0, 1, 1, 1, 2, 2, 2, 0, 1)
sync_reset;
check_mem(1029,"011100010","000011100",0,'1'); -- (0, 1, 1, 1, 2, 2, 2, 1, 0)
sync_reset;
check_mem(1030,"011100010","000011101",0,'1'); -- (0, 1, 1, 1, 2, 2, 2, 1, 2)
sync_reset;
check_mem(1031,"011100001","000011110",0,'1'); -- (0, 1, 1, 1, 2, 2, 2, 2, 1)
sync_reset;
check_mem(1032,"011000000","000100000",0,'1'); -- (0, 1, 1, 2, 0, 0, 0, 0, 0)
sync_reset;
check_mem(1033,"011000000","000100001",0,'1'); -- (0, 1, 1, 2, 0, 0, 0, 0, 2)
sync_reset;
check_mem(1034,"011000010","000100001",0,'1'); -- (0, 1, 1, 2, 0, 0, 0, 1, 2)
sync_reset;
check_mem(1035,"011000000","000100010",0,'1'); -- (0, 1, 1, 2, 0, 0, 0, 2, 0)
sync_reset;
check_mem(1036,"011000001","000100010",0,'1'); -- (0, 1, 1, 2, 0, 0, 0, 2, 1)
sync_reset;
check_mem(1037,"011000100","000100001",0,'1'); -- (0, 1, 1, 2, 0, 0, 1, 0, 2)
sync_reset;
check_mem(1038,"011000100","000100010",0,'1'); -- (0, 1, 1, 2, 0, 0, 1, 2, 0)
sync_reset;
check_mem(1039,"011000100","000100011",0,'1'); -- (0, 1, 1, 2, 0, 0, 1, 2, 2)
sync_reset;
check_mem(1040,"011000000","000100100",0,'1'); -- (0, 1, 1, 2, 0, 0, 2, 0, 0)
sync_reset;
check_mem(1041,"011000001","000100100",0,'1'); -- (0, 1, 1, 2, 0, 0, 2, 0, 1)
sync_reset;
check_mem(1042,"011000010","000100100",0,'1'); -- (0, 1, 1, 2, 0, 0, 2, 1, 0)
sync_reset;
check_mem(1043,"011000010","000100101",0,'1'); -- (0, 1, 1, 2, 0, 0, 2, 1, 2)
sync_reset;
check_mem(1044,"011000001","000100110",0,'1'); -- (0, 1, 1, 2, 0, 0, 2, 2, 1)
sync_reset;
check_mem(1045,"011001000","000100001",0,'1'); -- (0, 1, 1, 2, 0, 1, 0, 0, 2)
sync_reset;
check_mem(1046,"011001000","000100010",0,'1'); -- (0, 1, 1, 2, 0, 1, 0, 2, 0)
sync_reset;
check_mem(1047,"011001000","000100011",0,'1'); -- (0, 1, 1, 2, 0, 1, 0, 2, 2)
sync_reset;
check_mem(1048,"011001100","000100011",0,'1'); -- (0, 1, 1, 2, 0, 1, 1, 2, 2)
sync_reset;
check_mem(1049,"011001000","000100100",0,'1'); -- (0, 1, 1, 2, 0, 1, 2, 0, 0)
sync_reset;
check_mem(1050,"011001000","000100101",0,'1'); -- (0, 1, 1, 2, 0, 1, 2, 0, 2)
sync_reset;
check_mem(1051,"011001010","000100101",0,'1'); -- (0, 1, 1, 2, 0, 1, 2, 1, 2)
sync_reset;
check_mem(1052,"011001000","000100110",0,'1'); -- (0, 1, 1, 2, 0, 1, 2, 2, 0)
sync_reset;
check_mem(1053,"011000000","000101000",0,'1'); -- (0, 1, 1, 2, 0, 2, 0, 0, 0)
sync_reset;
check_mem(1054,"011000001","000101000",0,'1'); -- (0, 1, 1, 2, 0, 2, 0, 0, 1)
sync_reset;
check_mem(1055,"011000010","000101000",4,'1'); -- (0, 1, 1, 2, 0, 2, 0, 1, 0)
sync_reset;
check_mem(1056,"011000010","000101001",0,'1'); -- (0, 1, 1, 2, 0, 2, 0, 1, 2)
sync_reset;
check_mem(1057,"011000001","000101010",0,'1'); -- (0, 1, 1, 2, 0, 2, 0, 2, 1)
sync_reset;
check_mem(1058,"011000100","000101000",4,'1'); -- (0, 1, 1, 2, 0, 2, 1, 0, 0)
sync_reset;
check_mem(1059,"011000100","000101001",0,'1'); -- (0, 1, 1, 2, 0, 2, 1, 0, 2)
sync_reset;
check_mem(1060,"011000110","000101001",4,'1'); -- (0, 1, 1, 2, 0, 2, 1, 1, 2)
sync_reset;
check_mem(1061,"011000100","000101010",0,'1'); -- (0, 1, 1, 2, 0, 2, 1, 2, 0)
sync_reset;
check_mem(1062,"011000101","000101010",4,'1'); -- (0, 1, 1, 2, 0, 2, 1, 2, 1)
sync_reset;
check_mem(1063,"011000001","000101100",0,'1'); -- (0, 1, 1, 2, 0, 2, 2, 0, 1)
sync_reset;
check_mem(1064,"011000010","000101100",0,'1'); -- (0, 1, 1, 2, 0, 2, 2, 1, 0)
sync_reset;
check_mem(1065,"011000011","000101100",0,'1'); -- (0, 1, 1, 2, 0, 2, 2, 1, 1)
sync_reset;
check_mem(1066,"011010000","000100001",0,'1'); -- (0, 1, 1, 2, 1, 0, 0, 0, 2)
sync_reset;
check_mem(1067,"011010000","000100010",0,'1'); -- (0, 1, 1, 2, 1, 0, 0, 2, 0)
sync_reset;
check_mem(1068,"011010000","000100011",0,'1'); -- (0, 1, 1, 2, 1, 0, 0, 2, 2)
sync_reset;
check_mem(1069,"011010000","000100100",0,'1'); -- (0, 1, 1, 2, 1, 0, 2, 0, 0)
sync_reset;
check_mem(1070,"011010000","000100101",0,'1'); -- (0, 1, 1, 2, 1, 0, 2, 0, 2)
sync_reset;
check_mem(1071,"011010000","000100110",0,'1'); -- (0, 1, 1, 2, 1, 0, 2, 2, 0)
sync_reset;
check_mem(1072,"011010001","000100110",0,'1'); -- (0, 1, 1, 2, 1, 0, 2, 2, 1)
sync_reset;
check_mem(1073,"011011000","000100011",6,'1'); -- (0, 1, 1, 2, 1, 1, 0, 2, 2)
sync_reset;
check_mem(1074,"011011000","000100101",0,'1'); -- (0, 1, 1, 2, 1, 1, 2, 0, 2)
sync_reset;
check_mem(1075,"011011000","000100110",0,'1'); -- (0, 1, 1, 2, 1, 1, 2, 2, 0)
sync_reset;
check_mem(1076,"011010000","000101000",0,'1'); -- (0, 1, 1, 2, 1, 2, 0, 0, 0)
sync_reset;
check_mem(1077,"011010000","000101001",0,'1'); -- (0, 1, 1, 2, 1, 2, 0, 0, 2)
sync_reset;
check_mem(1078,"011010000","000101010",0,'1'); -- (0, 1, 1, 2, 1, 2, 0, 2, 0)
sync_reset;
check_mem(1079,"011010001","000101010",0,'1'); -- (0, 1, 1, 2, 1, 2, 0, 2, 1)
sync_reset;
check_mem(1080,"011010000","000101100",0,'1'); -- (0, 1, 1, 2, 1, 2, 2, 0, 0)
sync_reset;
check_mem(1081,"011010001","000101100",0,'1'); -- (0, 1, 1, 2, 1, 2, 2, 0, 1)
sync_reset;
check_mem(1082,"011010001","000101110",0,'1'); -- (0, 1, 1, 2, 1, 2, 2, 2, 1)
sync_reset;
check_mem(1083,"011000000","000110000",0,'1'); -- (0, 1, 1, 2, 2, 0, 0, 0, 0)
sync_reset;
check_mem(1084,"011000001","000110000",5,'1'); -- (0, 1, 1, 2, 2, 0, 0, 0, 1)
sync_reset;
check_mem(1085,"011000010","000110000",0,'1'); -- (0, 1, 1, 2, 2, 0, 0, 1, 0)
sync_reset;
check_mem(1086,"011000010","000110001",0,'1'); -- (0, 1, 1, 2, 2, 0, 0, 1, 2)
sync_reset;
check_mem(1087,"011000001","000110010",0,'1'); -- (0, 1, 1, 2, 2, 0, 0, 2, 1)
sync_reset;
check_mem(1088,"011000100","000110000",0,'1'); -- (0, 1, 1, 2, 2, 0, 1, 0, 0)
sync_reset;
check_mem(1089,"011000100","000110001",0,'1'); -- (0, 1, 1, 2, 2, 0, 1, 0, 2)
sync_reset;
check_mem(1090,"011000110","000110001",0,'1'); -- (0, 1, 1, 2, 2, 0, 1, 1, 2)
sync_reset;
check_mem(1091,"011000100","000110010",0,'1'); -- (0, 1, 1, 2, 2, 0, 1, 2, 0)
sync_reset;
check_mem(1092,"011000101","000110010",5,'1'); -- (0, 1, 1, 2, 2, 0, 1, 2, 1)
sync_reset;
check_mem(1093,"011000001","000110100",0,'1'); -- (0, 1, 1, 2, 2, 0, 2, 0, 1)
sync_reset;
check_mem(1094,"011000010","000110100",0,'1'); -- (0, 1, 1, 2, 2, 0, 2, 1, 0)
sync_reset;
check_mem(1095,"011000011","000110100",0,'1'); -- (0, 1, 1, 2, 2, 0, 2, 1, 1)
sync_reset;
check_mem(1096,"011001000","000110000",0,'1'); -- (0, 1, 1, 2, 2, 1, 0, 0, 0)
sync_reset;
check_mem(1097,"011001000","000110001",0,'1'); -- (0, 1, 1, 2, 2, 1, 0, 0, 2)
sync_reset;
check_mem(1098,"011001010","000110001",0,'1'); -- (0, 1, 1, 2, 2, 1, 0, 1, 2)
sync_reset;
check_mem(1099,"011001000","000110010",0,'1'); -- (0, 1, 1, 2, 2, 1, 0, 2, 0)
sync_reset;
check_mem(1100,"011001100","000110001",0,'1'); -- (0, 1, 1, 2, 2, 1, 1, 0, 2)
sync_reset;
check_mem(1101,"011001100","000110010",0,'1'); -- (0, 1, 1, 2, 2, 1, 1, 2, 0)
sync_reset;
check_mem(1102,"011001100","000110011",0,'1'); -- (0, 1, 1, 2, 2, 1, 1, 2, 2)
sync_reset;
check_mem(1103,"011001000","000110100",0,'1'); -- (0, 1, 1, 2, 2, 1, 2, 0, 0)
sync_reset;
check_mem(1104,"011001010","000110100",0,'1'); -- (0, 1, 1, 2, 2, 1, 2, 1, 0)
sync_reset;
check_mem(1105,"011001010","000110101",0,'1'); -- (0, 1, 1, 2, 2, 1, 2, 1, 2)
sync_reset;
check_mem(1106,"010000000","001000000",4,'1'); -- (0, 1, 2, 0, 0, 0, 0, 0, 0)
sync_reset;
check_mem(1107,"010000001","001000000",4,'1'); -- (0, 1, 2, 0, 0, 0, 0, 0, 1)
sync_reset;
check_mem(1108,"010000010","001000000",4,'1'); -- (0, 1, 2, 0, 0, 0, 0, 1, 0)
sync_reset;
check_mem(1109,"010000010","001000001",4,'1'); -- (0, 1, 2, 0, 0, 0, 0, 1, 2)
sync_reset;
check_mem(1110,"010000001","001000010",0,'1'); -- (0, 1, 2, 0, 0, 0, 0, 2, 1)
sync_reset;
check_mem(1111,"010000100","001000000",4,'1'); -- (0, 1, 2, 0, 0, 0, 1, 0, 0)
sync_reset;
check_mem(1112,"010000100","001000001",5,'1'); -- (0, 1, 2, 0, 0, 0, 1, 0, 2)
sync_reset;
check_mem(1113,"010000110","001000001",4,'1'); -- (0, 1, 2, 0, 0, 0, 1, 1, 2)
sync_reset;
check_mem(1114,"010000100","001000010",0,'1'); -- (0, 1, 2, 0, 0, 0, 1, 2, 0)
sync_reset;
check_mem(1115,"010000101","001000010",0,'1'); -- (0, 1, 2, 0, 0, 0, 1, 2, 1)
sync_reset;
check_mem(1116,"010000001","001000100",4,'1'); -- (0, 1, 2, 0, 0, 0, 2, 0, 1)
sync_reset;
check_mem(1117,"010000010","001000100",4,'1'); -- (0, 1, 2, 0, 0, 0, 2, 1, 0)
sync_reset;
check_mem(1118,"010000011","001000100",4,'1'); -- (0, 1, 2, 0, 0, 0, 2, 1, 1)
sync_reset;
check_mem(1119,"010001000","001000000",3,'1'); -- (0, 1, 2, 0, 0, 1, 0, 0, 0)
sync_reset;
check_mem(1120,"010001000","001000001",4,'1'); -- (0, 1, 2, 0, 0, 1, 0, 0, 2)
sync_reset;
check_mem(1121,"010001010","001000001",4,'1'); -- (0, 1, 2, 0, 0, 1, 0, 1, 2)
sync_reset;
check_mem(1122,"010001000","001000010",3,'1'); -- (0, 1, 2, 0, 0, 1, 0, 2, 0)
sync_reset;
check_mem(1123,"010001001","001000010",0,'1'); -- (0, 1, 2, 0, 0, 1, 0, 2, 1)
sync_reset;
check_mem(1124,"010001100","001000001",3,'1'); -- (0, 1, 2, 0, 0, 1, 1, 0, 2)
sync_reset;
check_mem(1125,"010001100","001000010",0,'1'); -- (0, 1, 2, 0, 0, 1, 1, 2, 0)
sync_reset;
check_mem(1126,"010001100","001000011",3,'1'); -- (0, 1, 2, 0, 0, 1, 1, 2, 2)
sync_reset;
check_mem(1127,"010001000","001000100",4,'1'); -- (0, 1, 2, 0, 0, 1, 2, 0, 0)
sync_reset;
check_mem(1128,"010001001","001000100",0,'1'); -- (0, 1, 2, 0, 0, 1, 2, 0, 1)
sync_reset;
check_mem(1129,"010001010","001000100",4,'1'); -- (0, 1, 2, 0, 0, 1, 2, 1, 0)
sync_reset;
check_mem(1130,"010001010","001000101",4,'1'); -- (0, 1, 2, 0, 0, 1, 2, 1, 2)
sync_reset;
check_mem(1131,"010001001","001000110",4,'1'); -- (0, 1, 2, 0, 0, 1, 2, 2, 1)
sync_reset;
check_mem(1132,"010000001","001001000",3,'1'); -- (0, 1, 2, 0, 0, 2, 0, 0, 1)
sync_reset;
check_mem(1133,"010000010","001001000",4,'1'); -- (0, 1, 2, 0, 0, 2, 0, 1, 0)
sync_reset;
check_mem(1134,"010000011","001001000",0,'1'); -- (0, 1, 2, 0, 0, 2, 0, 1, 1)
sync_reset;
check_mem(1135,"010000100","001001000",8,'1'); -- (0, 1, 2, 0, 0, 2, 1, 0, 0)
sync_reset;
check_mem(1136,"010000101","001001000",0,'1'); -- (0, 1, 2, 0, 0, 2, 1, 0, 1)
sync_reset;
check_mem(1137,"010000110","001001000",8,'1'); -- (0, 1, 2, 0, 0, 2, 1, 1, 0)
sync_reset;
check_mem(1138,"010000101","001001010",0,'1'); -- (0, 1, 2, 0, 0, 2, 1, 2, 1)
sync_reset;
check_mem(1139,"010000011","001001100",4,'1'); -- (0, 1, 2, 0, 0, 2, 2, 1, 1)
sync_reset;
check_mem(1140,"010010000","001000000",7,'1'); -- (0, 1, 2, 0, 1, 0, 0, 0, 0)
sync_reset;
check_mem(1141,"010010000","001000001",5,'1'); -- (0, 1, 2, 0, 1, 0, 0, 0, 2)
sync_reset;
check_mem(1142,"010010000","001000010",3,'1'); -- (0, 1, 2, 0, 1, 0, 0, 2, 0)
sync_reset;
check_mem(1143,"010010001","001000010",0,'1'); -- (0, 1, 2, 0, 1, 0, 0, 2, 1)
sync_reset;
check_mem(1144,"010010100","001000001",5,'1'); -- (0, 1, 2, 0, 1, 0, 1, 0, 2)
sync_reset;
check_mem(1145,"010010100","001000010",0,'1'); -- (0, 1, 2, 0, 1, 0, 1, 2, 0)
sync_reset;
check_mem(1146,"010010100","001000011",5,'1'); -- (0, 1, 2, 0, 1, 0, 1, 2, 2)
sync_reset;
check_mem(1147,"010010000","001000100",0,'1'); -- (0, 1, 2, 0, 1, 0, 2, 0, 0)
sync_reset;
check_mem(1148,"010010001","001000100",0,'1'); -- (0, 1, 2, 0, 1, 0, 2, 0, 1)
sync_reset;
check_mem(1149,"010010001","001000110",0,'1'); -- (0, 1, 2, 0, 1, 0, 2, 2, 1)
sync_reset;
check_mem(1150,"010011000","001000001",0,'1'); -- (0, 1, 2, 0, 1, 1, 0, 0, 2)
sync_reset;
check_mem(1151,"010011000","001000010",3,'1'); -- (0, 1, 2, 0, 1, 1, 0, 2, 0)
sync_reset;
check_mem(1152,"010011000","001000011",3,'1'); -- (0, 1, 2, 0, 1, 1, 0, 2, 2)
sync_reset;
check_mem(1153,"010011100","001000011",3,'1'); -- (0, 1, 2, 0, 1, 1, 1, 2, 2)
sync_reset;
check_mem(1154,"010011000","001000100",0,'1'); -- (0, 1, 2, 0, 1, 1, 2, 0, 0)
sync_reset;
check_mem(1155,"010011000","001000101",3,'1'); -- (0, 1, 2, 0, 1, 1, 2, 0, 2)
sync_reset;
check_mem(1156,"010011000","001000110",3,'1'); -- (0, 1, 2, 0, 1, 1, 2, 2, 0)
sync_reset;
check_mem(1157,"010011001","001000110",0,'1'); -- (0, 1, 2, 0, 1, 1, 2, 2, 1)
sync_reset;
check_mem(1158,"010010000","001001000",7,'1'); -- (0, 1, 2, 0, 1, 2, 0, 0, 0)
sync_reset;
check_mem(1159,"010010001","001001000",0,'1'); -- (0, 1, 2, 0, 1, 2, 0, 0, 1)
sync_reset;
check_mem(1160,"010010001","001001010",0,'1'); -- (0, 1, 2, 0, 1, 2, 0, 2, 1)
sync_reset;
check_mem(1161,"010010100","001001000",8,'1'); -- (0, 1, 2, 0, 1, 2, 1, 0, 0)
sync_reset;
check_mem(1162,"010010100","001001010",8,'1'); -- (0, 1, 2, 0, 1, 2, 1, 2, 0)
sync_reset;
check_mem(1163,"010010101","001001010",0,'1'); -- (0, 1, 2, 0, 1, 2, 1, 2, 1)
sync_reset;
check_mem(1164,"010010001","001001100",0,'1'); -- (0, 1, 2, 0, 1, 2, 2, 0, 1)
sync_reset;
check_mem(1165,"010000001","001010000",6,'1'); -- (0, 1, 2, 0, 2, 0, 0, 0, 1)
sync_reset;
check_mem(1166,"010000010","001010000",0,'1'); -- (0, 1, 2, 0, 2, 0, 0, 1, 0)
sync_reset;
check_mem(1167,"010000011","001010000",6,'1'); -- (0, 1, 2, 0, 2, 0, 0, 1, 1)
sync_reset;
check_mem(1168,"010000100","001010000",0,'1'); -- (0, 1, 2, 0, 2, 0, 1, 0, 0)
sync_reset;
check_mem(1169,"010000101","001010000",7,'1'); -- (0, 1, 2, 0, 2, 0, 1, 0, 1)
sync_reset;
check_mem(1170,"010000110","001010000",8,'1'); -- (0, 1, 2, 0, 2, 0, 1, 1, 0)
sync_reset;
check_mem(1171,"010000110","001010001",0,'1'); -- (0, 1, 2, 0, 2, 0, 1, 1, 2)
sync_reset;
check_mem(1172,"010000101","001010010",0,'1'); -- (0, 1, 2, 0, 2, 0, 1, 2, 1)
sync_reset;
check_mem(1173,"010001000","001010000",6,'1'); -- (0, 1, 2, 0, 2, 1, 0, 0, 0)
sync_reset;
check_mem(1174,"010001001","001010000",6,'1'); -- (0, 1, 2, 0, 2, 1, 0, 0, 1)
sync_reset;
check_mem(1175,"010001010","001010000",0,'1'); -- (0, 1, 2, 0, 2, 1, 0, 1, 0)
sync_reset;
check_mem(1176,"010001010","001010001",0,'1'); -- (0, 1, 2, 0, 2, 1, 0, 1, 2)
sync_reset;
check_mem(1177,"010001001","001010010",6,'1'); -- (0, 1, 2, 0, 2, 1, 0, 2, 1)
sync_reset;
check_mem(1178,"010001100","001010000",0,'1'); -- (0, 1, 2, 0, 2, 1, 1, 0, 0)
sync_reset;
check_mem(1179,"010001100","001010001",0,'1'); -- (0, 1, 2, 0, 2, 1, 1, 0, 2)
sync_reset;
check_mem(1180,"010001110","001010001",0,'1'); -- (0, 1, 2, 0, 2, 1, 1, 1, 2)
sync_reset;
check_mem(1181,"010001100","001010010",0,'1'); -- (0, 1, 2, 0, 2, 1, 1, 2, 0)
sync_reset;
check_mem(1182,"010001101","001010010",0,'1'); -- (0, 1, 2, 0, 2, 1, 1, 2, 1)
sync_reset;
check_mem(1183,"010000011","001011000",6,'1'); -- (0, 1, 2, 0, 2, 2, 0, 1, 1)
sync_reset;
check_mem(1184,"010000101","001011000",3,'1'); -- (0, 1, 2, 0, 2, 2, 1, 0, 1)
sync_reset;
check_mem(1185,"010000110","001011000",8,'1'); -- (0, 1, 2, 0, 2, 2, 1, 1, 0)
sync_reset;
check_mem(1186,"010100000","001000000",8,'1'); -- (0, 1, 2, 1, 0, 0, 0, 0, 0)
sync_reset;
check_mem(1187,"010100000","001000001",0,'1'); -- (0, 1, 2, 1, 0, 0, 0, 0, 2)
sync_reset;
check_mem(1188,"010100010","001000001",4,'1'); -- (0, 1, 2, 1, 0, 0, 0, 1, 2)
sync_reset;
check_mem(1189,"010100000","001000010",4,'1'); -- (0, 1, 2, 1, 0, 0, 0, 2, 0)
sync_reset;
check_mem(1190,"010100001","001000010",0,'1'); -- (0, 1, 2, 1, 0, 0, 0, 2, 1)
sync_reset;
check_mem(1191,"010100100","001000001",0,'1'); -- (0, 1, 2, 1, 0, 0, 1, 0, 2)
sync_reset;
check_mem(1192,"010100100","001000010",0,'1'); -- (0, 1, 2, 1, 0, 0, 1, 2, 0)
sync_reset;
check_mem(1193,"010100100","001000011",0,'1'); -- (0, 1, 2, 1, 0, 0, 1, 2, 2)
sync_reset;
check_mem(1194,"010100000","001000100",4,'1'); -- (0, 1, 2, 1, 0, 0, 2, 0, 0)
sync_reset;
check_mem(1195,"010100001","001000100",4,'1'); -- (0, 1, 2, 1, 0, 0, 2, 0, 1)
sync_reset;
check_mem(1196,"010100010","001000100",4,'1'); -- (0, 1, 2, 1, 0, 0, 2, 1, 0)
sync_reset;
check_mem(1197,"010100010","001000101",4,'1'); -- (0, 1, 2, 1, 0, 0, 2, 1, 2)
sync_reset;
check_mem(1198,"010100001","001000110",4,'1'); -- (0, 1, 2, 1, 0, 0, 2, 2, 1)
sync_reset;
check_mem(1199,"010101000","001000001",4,'1'); -- (0, 1, 2, 1, 0, 1, 0, 0, 2)
sync_reset;
check_mem(1200,"010101000","001000010",4,'1'); -- (0, 1, 2, 1, 0, 1, 0, 2, 0)
sync_reset;
check_mem(1201,"010101000","001000011",4,'1'); -- (0, 1, 2, 1, 0, 1, 0, 2, 2)
sync_reset;
check_mem(1202,"010101100","001000011",0,'1'); -- (0, 1, 2, 1, 0, 1, 1, 2, 2)
sync_reset;
check_mem(1203,"010101000","001000100",4,'1'); -- (0, 1, 2, 1, 0, 1, 2, 0, 0)
sync_reset;
check_mem(1204,"010101000","001000101",4,'1'); -- (0, 1, 2, 1, 0, 1, 2, 0, 2)
sync_reset;
check_mem(1205,"010101010","001000101",4,'1'); -- (0, 1, 2, 1, 0, 1, 2, 1, 2)
sync_reset;
check_mem(1206,"010101000","001000110",4,'1'); -- (0, 1, 2, 1, 0, 1, 2, 2, 0)
sync_reset;
check_mem(1207,"010101001","001000110",4,'1'); -- (0, 1, 2, 1, 0, 1, 2, 2, 1)
sync_reset;
check_mem(1208,"010100000","001001000",8,'1'); -- (0, 1, 2, 1, 0, 2, 0, 0, 0)
sync_reset;
check_mem(1209,"010100001","001001000",0,'1'); -- (0, 1, 2, 1, 0, 2, 0, 0, 1)
sync_reset;
check_mem(1210,"010100010","001001000",4,'1'); -- (0, 1, 2, 1, 0, 2, 0, 1, 0)
sync_reset;
check_mem(1211,"010100001","001001010",0,'1'); -- (0, 1, 2, 1, 0, 2, 0, 2, 1)
sync_reset;
check_mem(1212,"010100100","001001000",8,'1'); -- (0, 1, 2, 1, 0, 2, 1, 0, 0)
sync_reset;
check_mem(1213,"010100100","001001010",0,'1'); -- (0, 1, 2, 1, 0, 2, 1, 2, 0)
sync_reset;
check_mem(1214,"010100101","001001010",0,'1'); -- (0, 1, 2, 1, 0, 2, 1, 2, 1)
sync_reset;
check_mem(1215,"010100001","001001100",4,'1'); -- (0, 1, 2, 1, 0, 2, 2, 0, 1)
sync_reset;
check_mem(1216,"010100010","001001100",4,'1'); -- (0, 1, 2, 1, 0, 2, 2, 1, 0)
sync_reset;
check_mem(1217,"010100011","001001100",4,'1'); -- (0, 1, 2, 1, 0, 2, 2, 1, 1)
sync_reset;
check_mem(1218,"010110000","001000001",5,'1'); -- (0, 1, 2, 1, 1, 0, 0, 0, 2)
sync_reset;
check_mem(1219,"010110000","001000010",5,'1'); -- (0, 1, 2, 1, 1, 0, 0, 2, 0)
sync_reset;
check_mem(1220,"010110000","001000011",5,'1'); -- (0, 1, 2, 1, 1, 0, 0, 2, 2)
sync_reset;
check_mem(1221,"010110100","001000011",5,'1'); -- (0, 1, 2, 1, 1, 0, 1, 2, 2)
sync_reset;
check_mem(1222,"010110000","001000100",0,'1'); -- (0, 1, 2, 1, 1, 0, 2, 0, 0)
sync_reset;
check_mem(1223,"010110000","001000101",5,'1'); -- (0, 1, 2, 1, 1, 0, 2, 0, 2)
sync_reset;
check_mem(1224,"010110000","001000110",5,'1'); -- (0, 1, 2, 1, 1, 0, 2, 2, 0)
sync_reset;
check_mem(1225,"010110001","001000110",0,'1'); -- (0, 1, 2, 1, 1, 0, 2, 2, 1)
sync_reset;
check_mem(1226,"010110000","001001000",8,'1'); -- (0, 1, 2, 1, 1, 2, 0, 0, 0)
sync_reset;
check_mem(1227,"010110000","001001010",8,'1'); -- (0, 1, 2, 1, 1, 2, 0, 2, 0)
sync_reset;
check_mem(1228,"010110001","001001010",0,'1'); -- (0, 1, 2, 1, 1, 2, 0, 2, 1)
sync_reset;
check_mem(1229,"010110100","001001010",8,'1'); -- (0, 1, 2, 1, 1, 2, 1, 2, 0)
sync_reset;
check_mem(1230,"010110000","001001100",7,'1'); -- (0, 1, 2, 1, 1, 2, 2, 0, 0)
sync_reset;
check_mem(1231,"010110001","001001100",0,'1'); -- (0, 1, 2, 1, 1, 2, 2, 0, 1)
sync_reset;
check_mem(1232,"010110001","001001110",0,'1'); -- (0, 1, 2, 1, 1, 2, 2, 2, 1)
sync_reset;
check_mem(1233,"010100000","001010000",6,'1'); -- (0, 1, 2, 1, 2, 0, 0, 0, 0)
sync_reset;
check_mem(1234,"010100001","001010000",6,'1'); -- (0, 1, 2, 1, 2, 0, 0, 0, 1)
sync_reset;
check_mem(1235,"010100010","001010000",0,'1'); -- (0, 1, 2, 1, 2, 0, 0, 1, 0)
sync_reset;
check_mem(1236,"010100010","001010001",0,'1'); -- (0, 1, 2, 1, 2, 0, 0, 1, 2)
sync_reset;
check_mem(1237,"010100001","001010010",6,'1'); -- (0, 1, 2, 1, 2, 0, 0, 2, 1)
sync_reset;
check_mem(1238,"010100100","001010000",0,'1'); -- (0, 1, 2, 1, 2, 0, 1, 0, 0)
sync_reset;
check_mem(1239,"010100100","001010001",0,'1'); -- (0, 1, 2, 1, 2, 0, 1, 0, 2)
sync_reset;
check_mem(1240,"010100110","001010001",0,'1'); -- (0, 1, 2, 1, 2, 0, 1, 1, 2)
sync_reset;
check_mem(1241,"010100100","001010010",0,'1'); -- (0, 1, 2, 1, 2, 0, 1, 2, 0)
sync_reset;
check_mem(1242,"010100101","001010010",0,'1'); -- (0, 1, 2, 1, 2, 0, 1, 2, 1)
sync_reset;
check_mem(1243,"010101000","001010000",0,'1'); -- (0, 1, 2, 1, 2, 1, 0, 0, 0)
sync_reset;
check_mem(1244,"010101000","001010001",0,'1'); -- (0, 1, 2, 1, 2, 1, 0, 0, 2)
sync_reset;
check_mem(1245,"010101010","001010001",0,'1'); -- (0, 1, 2, 1, 2, 1, 0, 1, 2)
sync_reset;
check_mem(1246,"010101000","001010010",6,'1'); -- (0, 1, 2, 1, 2, 1, 0, 2, 0)
sync_reset;
check_mem(1247,"010101001","001010010",6,'1'); -- (0, 1, 2, 1, 2, 1, 0, 2, 1)
sync_reset;
check_mem(1248,"010101100","001010001",0,'1'); -- (0, 1, 2, 1, 2, 1, 1, 0, 2)
sync_reset;
check_mem(1249,"010101100","001010010",0,'1'); -- (0, 1, 2, 1, 2, 1, 1, 2, 0)
sync_reset;
check_mem(1250,"010101100","001010011",0,'1'); -- (0, 1, 2, 1, 2, 1, 1, 2, 2)
sync_reset;
check_mem(1251,"010100001","001011000",6,'1'); -- (0, 1, 2, 1, 2, 2, 0, 0, 1)
sync_reset;
check_mem(1252,"010100010","001011000",0,'1'); -- (0, 1, 2, 1, 2, 2, 0, 1, 0)
sync_reset;
check_mem(1253,"010100011","001011000",6,'1'); -- (0, 1, 2, 1, 2, 2, 0, 1, 1)
sync_reset;
check_mem(1254,"010100100","001011000",0,'1'); -- (0, 1, 2, 1, 2, 2, 1, 0, 0)
sync_reset;
check_mem(1255,"010100101","001011000",0,'1'); -- (0, 1, 2, 1, 2, 2, 1, 0, 1)
sync_reset;
check_mem(1256,"010100110","001011000",8,'1'); -- (0, 1, 2, 1, 2, 2, 1, 1, 0)
sync_reset;
check_mem(1257,"010100101","001011010",0,'1'); -- (0, 1, 2, 1, 2, 2, 1, 2, 1)
sync_reset;
check_mem(1258,"010000001","001100000",4,'1'); -- (0, 1, 2, 2, 0, 0, 0, 0, 1)
sync_reset;
check_mem(1259,"010000010","001100000",4,'1'); -- (0, 1, 2, 2, 0, 0, 0, 1, 0)
sync_reset;
check_mem(1260,"010000011","001100000",0,'1'); -- (0, 1, 2, 2, 0, 0, 0, 1, 1)
sync_reset;
check_mem(1261,"010000100","001100000",7,'1'); -- (0, 1, 2, 2, 0, 0, 1, 0, 0)
sync_reset;
check_mem(1262,"010000101","001100000",7,'1'); -- (0, 1, 2, 2, 0, 0, 1, 0, 1)
sync_reset;
check_mem(1263,"010000110","001100000",0,'1'); -- (0, 1, 2, 2, 0, 0, 1, 1, 0)
sync_reset;
check_mem(1264,"010000110","001100001",4,'1'); -- (0, 1, 2, 2, 0, 0, 1, 1, 2)
sync_reset;
check_mem(1265,"010000101","001100010",0,'1'); -- (0, 1, 2, 2, 0, 0, 1, 2, 1)
sync_reset;
check_mem(1266,"010000011","001100100",4,'1'); -- (0, 1, 2, 2, 0, 0, 2, 1, 1)
sync_reset;
check_mem(1267,"010001000","001100000",0,'1'); -- (0, 1, 2, 2, 0, 1, 0, 0, 0)
sync_reset;
check_mem(1268,"010001001","001100000",6,'1'); -- (0, 1, 2, 2, 0, 1, 0, 0, 1)
sync_reset;
check_mem(1269,"010001010","001100000",4,'1'); -- (0, 1, 2, 2, 0, 1, 0, 1, 0)
sync_reset;
check_mem(1270,"010001010","001100001",4,'1'); -- (0, 1, 2, 2, 0, 1, 0, 1, 2)
sync_reset;
check_mem(1271,"010001001","001100010",0,'1'); -- (0, 1, 2, 2, 0, 1, 0, 2, 1)
sync_reset;
check_mem(1272,"010001100","001100000",4,'1'); -- (0, 1, 2, 2, 0, 1, 1, 0, 0)
sync_reset;
check_mem(1273,"010001100","001100001",0,'1'); -- (0, 1, 2, 2, 0, 1, 1, 0, 2)
sync_reset;
check_mem(1274,"010001110","001100001",4,'1'); -- (0, 1, 2, 2, 0, 1, 1, 1, 2)
sync_reset;
check_mem(1275,"010001100","001100010",0,'1'); -- (0, 1, 2, 2, 0, 1, 1, 2, 0)
sync_reset;
check_mem(1276,"010001101","001100010",0,'1'); -- (0, 1, 2, 2, 0, 1, 1, 2, 1)
sync_reset;
check_mem(1277,"010001001","001100100",0,'1'); -- (0, 1, 2, 2, 0, 1, 2, 0, 1)
sync_reset;
check_mem(1278,"010001010","001100100",4,'1'); -- (0, 1, 2, 2, 0, 1, 2, 1, 0)
sync_reset;
check_mem(1279,"010001011","001100100",0,'1'); -- (0, 1, 2, 2, 0, 1, 2, 1, 1)
sync_reset;
check_mem(1280,"010000011","001101000",4,'1'); -- (0, 1, 2, 2, 0, 2, 0, 1, 1)
sync_reset;
check_mem(1281,"010000101","001101000",4,'1'); -- (0, 1, 2, 2, 0, 2, 1, 0, 1)
sync_reset;
check_mem(1282,"010000110","001101000",4,'1'); -- (0, 1, 2, 2, 0, 2, 1, 1, 0)
sync_reset;
check_mem(1283,"010010000","001100000",0,'1'); -- (0, 1, 2, 2, 1, 0, 0, 0, 0)
sync_reset;
check_mem(1284,"010010001","001100000",0,'1'); -- (0, 1, 2, 2, 1, 0, 0, 0, 1)
sync_reset;
check_mem(1285,"010010001","001100010",0,'1'); -- (0, 1, 2, 2, 1, 0, 0, 2, 1)
sync_reset;
check_mem(1286,"010010100","001100000",7,'1'); -- (0, 1, 2, 2, 1, 0, 1, 0, 0)
sync_reset;
check_mem(1287,"010010100","001100001",7,'1'); -- (0, 1, 2, 2, 1, 0, 1, 0, 2)
sync_reset;
check_mem(1288,"010010100","001100010",0,'1'); -- (0, 1, 2, 2, 1, 0, 1, 2, 0)
sync_reset;
check_mem(1289,"010010101","001100010",0,'1'); -- (0, 1, 2, 2, 1, 0, 1, 2, 1)
sync_reset;
check_mem(1290,"010010001","001100100",0,'1'); -- (0, 1, 2, 2, 1, 0, 2, 0, 1)
sync_reset;
check_mem(1291,"010011000","001100000",7,'1'); -- (0, 1, 2, 2, 1, 1, 0, 0, 0)
sync_reset;
check_mem(1292,"010011000","001100001",7,'1'); -- (0, 1, 2, 2, 1, 1, 0, 0, 2)
sync_reset;
check_mem(1293,"010011000","001100010",0,'1'); -- (0, 1, 2, 2, 1, 1, 0, 2, 0)
sync_reset;
check_mem(1294,"010011001","001100010",0,'1'); -- (0, 1, 2, 2, 1, 1, 0, 2, 1)
sync_reset;
check_mem(1295,"010011100","001100001",7,'1'); -- (0, 1, 2, 2, 1, 1, 1, 0, 2)
sync_reset;
check_mem(1296,"010011100","001100010",0,'1'); -- (0, 1, 2, 2, 1, 1, 1, 2, 0)
sync_reset;
check_mem(1297,"010011100","001100011",0,'1'); -- (0, 1, 2, 2, 1, 1, 1, 2, 2)
sync_reset;
check_mem(1298,"010011000","001100100",0,'1'); -- (0, 1, 2, 2, 1, 1, 2, 0, 0)
sync_reset;
check_mem(1299,"010011001","001100100",0,'1'); -- (0, 1, 2, 2, 1, 1, 2, 0, 1)
sync_reset;
check_mem(1300,"010011001","001100110",0,'1'); -- (0, 1, 2, 2, 1, 1, 2, 2, 1)
sync_reset;
check_mem(1301,"010010001","001101000",0,'1'); -- (0, 1, 2, 2, 1, 2, 0, 0, 1)
sync_reset;
check_mem(1302,"010010100","001101000",7,'1'); -- (0, 1, 2, 2, 1, 2, 1, 0, 0)
sync_reset;
check_mem(1303,"010010101","001101000",0,'1'); -- (0, 1, 2, 2, 1, 2, 1, 0, 1)
sync_reset;
check_mem(1304,"010010101","001101010",0,'1'); -- (0, 1, 2, 2, 1, 2, 1, 2, 1)
sync_reset;
check_mem(1305,"010000011","001110000",6,'1'); -- (0, 1, 2, 2, 2, 0, 0, 1, 1)
sync_reset;
check_mem(1306,"010000101","001110000",7,'1'); -- (0, 1, 2, 2, 2, 0, 1, 0, 1)
sync_reset;
check_mem(1307,"010000110","001110000",8,'1'); -- (0, 1, 2, 2, 2, 0, 1, 1, 0)
sync_reset;
check_mem(1308,"010001001","001110000",6,'1'); -- (0, 1, 2, 2, 2, 1, 0, 0, 1)
sync_reset;
check_mem(1309,"010001010","001110000",6,'1'); -- (0, 1, 2, 2, 2, 1, 0, 1, 0)
sync_reset;
check_mem(1310,"010001011","001110000",6,'1'); -- (0, 1, 2, 2, 2, 1, 0, 1, 1)
sync_reset;
check_mem(1311,"010001100","001110000",0,'1'); -- (0, 1, 2, 2, 2, 1, 1, 0, 0)
sync_reset;
check_mem(1312,"010001101","001110000",7,'1'); -- (0, 1, 2, 2, 2, 1, 1, 0, 1)
sync_reset;
check_mem(1313,"010001110","001110000",8,'1'); -- (0, 1, 2, 2, 2, 1, 1, 1, 0)
sync_reset;
check_mem(1314,"010001110","001110001",0,'1'); -- (0, 1, 2, 2, 2, 1, 1, 1, 2)
sync_reset;
check_mem(1315,"010001101","001110010",0,'1'); -- (0, 1, 2, 2, 2, 1, 1, 2, 1)
sync_reset;
check_mem(1316,"000000001","010000000",2,'1'); -- (0, 2, 0, 0, 0, 0, 0, 0, 1)
sync_reset;
check_mem(1317,"000000010","010000000",0,'1'); -- (0, 2, 0, 0, 0, 0, 0, 1, 0)
sync_reset;
check_mem(1318,"000000011","010000000",6,'1'); -- (0, 2, 0, 0, 0, 0, 0, 1, 1)
sync_reset;
check_mem(1319,"000000100","010000000",0,'1'); -- (0, 2, 0, 0, 0, 0, 1, 0, 0)
sync_reset;
check_mem(1320,"000000101","010000000",0,'1'); -- (0, 2, 0, 0, 0, 0, 1, 0, 1)
sync_reset;
check_mem(1321,"000000110","010000000",8,'1'); -- (0, 2, 0, 0, 0, 0, 1, 1, 0)
sync_reset;
check_mem(1322,"000000110","010000001",0,'1'); -- (0, 2, 0, 0, 0, 0, 1, 1, 2)
sync_reset;
check_mem(1323,"000000101","010000010",4,'1'); -- (0, 2, 0, 0, 0, 0, 1, 2, 1)
sync_reset;
check_mem(1324,"000000011","010000100",0,'1'); -- (0, 2, 0, 0, 0, 0, 2, 1, 1)
sync_reset;
check_mem(1325,"000001000","010000000",2,'1'); -- (0, 2, 0, 0, 0, 1, 0, 0, 0)
sync_reset;
check_mem(1326,"000001001","010000000",2,'1'); -- (0, 2, 0, 0, 0, 1, 0, 0, 1)
sync_reset;
check_mem(1327,"000001010","010000000",6,'1'); -- (0, 2, 0, 0, 0, 1, 0, 1, 0)
sync_reset;
check_mem(1328,"000001010","010000001",0,'1'); -- (0, 2, 0, 0, 0, 1, 0, 1, 2)
sync_reset;
check_mem(1329,"000001001","010000010",2,'1'); -- (0, 2, 0, 0, 0, 1, 0, 2, 1)
sync_reset;
check_mem(1330,"000001100","010000000",4,'1'); -- (0, 2, 0, 0, 0, 1, 1, 0, 0)
sync_reset;
check_mem(1331,"000001100","010000001",3,'1'); -- (0, 2, 0, 0, 0, 1, 1, 0, 2)
sync_reset;
check_mem(1332,"000001110","010000001",0,'1'); -- (0, 2, 0, 0, 0, 1, 1, 1, 2)
sync_reset;
check_mem(1333,"000001100","010000010",4,'1'); -- (0, 2, 0, 0, 0, 1, 1, 2, 0)
sync_reset;
check_mem(1334,"000001101","010000010",2,'1'); -- (0, 2, 0, 0, 0, 1, 1, 2, 1)
sync_reset;
check_mem(1335,"000001001","010000100",0,'1'); -- (0, 2, 0, 0, 0, 1, 2, 0, 1)
sync_reset;
check_mem(1336,"000001010","010000100",0,'1'); -- (0, 2, 0, 0, 0, 1, 2, 1, 0)
sync_reset;
check_mem(1337,"000001011","010000100",2,'1'); -- (0, 2, 0, 0, 0, 1, 2, 1, 1)
sync_reset;
check_mem(1338,"000000011","010001000",0,'1'); -- (0, 2, 0, 0, 0, 2, 0, 1, 1)
sync_reset;
check_mem(1339,"000000101","010001000",0,'1'); -- (0, 2, 0, 0, 0, 2, 1, 0, 1)
sync_reset;
check_mem(1340,"000000110","010001000",0,'1'); -- (0, 2, 0, 0, 0, 2, 1, 1, 0)
sync_reset;
check_mem(1341,"000010000","010000000",0,'1'); -- (0, 2, 0, 0, 1, 0, 0, 0, 0)
sync_reset;
check_mem(1342,"000010001","010000000",0,'1'); -- (0, 2, 0, 0, 1, 0, 0, 0, 1)
sync_reset;
check_mem(1343,"000010010","010000000",0,'1'); -- (0, 2, 0, 0, 1, 0, 0, 1, 0)
sync_reset;
check_mem(1344,"000010010","010000001",0,'1'); -- (0, 2, 0, 0, 1, 0, 0, 1, 2)
sync_reset;
check_mem(1345,"000010001","010000010",0,'1'); -- (0, 2, 0, 0, 1, 0, 0, 2, 1)
sync_reset;
check_mem(1346,"000010100","010000000",0,'1'); -- (0, 2, 0, 0, 1, 0, 1, 0, 0)
sync_reset;
check_mem(1347,"000010100","010000001",0,'1'); -- (0, 2, 0, 0, 1, 0, 1, 0, 2)
sync_reset;
check_mem(1348,"000010110","010000001",2,'1'); -- (0, 2, 0, 0, 1, 0, 1, 1, 2)
sync_reset;
check_mem(1349,"000010100","010000010",0,'1'); -- (0, 2, 0, 0, 1, 0, 1, 2, 0)
sync_reset;
check_mem(1350,"000010101","010000010",0,'1'); -- (0, 2, 0, 0, 1, 0, 1, 2, 1)
sync_reset;
check_mem(1351,"000010001","010000100",0,'1'); -- (0, 2, 0, 0, 1, 0, 2, 0, 1)
sync_reset;
check_mem(1352,"000010010","010000100",0,'1'); -- (0, 2, 0, 0, 1, 0, 2, 1, 0)
sync_reset;
check_mem(1353,"000010011","010000100",0,'1'); -- (0, 2, 0, 0, 1, 0, 2, 1, 1)
sync_reset;
check_mem(1354,"000011000","010000000",0,'1'); -- (0, 2, 0, 0, 1, 1, 0, 0, 0)
sync_reset;
check_mem(1355,"000011000","010000001",2,'1'); -- (0, 2, 0, 0, 1, 1, 0, 0, 2)
sync_reset;
check_mem(1356,"000011010","010000001",3,'1'); -- (0, 2, 0, 0, 1, 1, 0, 1, 2)
sync_reset;
check_mem(1357,"000011000","010000010",0,'1'); -- (0, 2, 0, 0, 1, 1, 0, 2, 0)
sync_reset;
check_mem(1358,"000011001","010000010",0,'1'); -- (0, 2, 0, 0, 1, 1, 0, 2, 1)
sync_reset;
check_mem(1359,"000011100","010000001",0,'1'); -- (0, 2, 0, 0, 1, 1, 1, 0, 2)
sync_reset;
check_mem(1360,"000011100","010000010",0,'1'); -- (0, 2, 0, 0, 1, 1, 1, 2, 0)
sync_reset;
check_mem(1361,"000011100","010000011",0,'1'); -- (0, 2, 0, 0, 1, 1, 1, 2, 2)
sync_reset;
check_mem(1362,"000011000","010000100",0,'1'); -- (0, 2, 0, 0, 1, 1, 2, 0, 0)
sync_reset;
check_mem(1363,"000011001","010000100",0,'1'); -- (0, 2, 0, 0, 1, 1, 2, 0, 1)
sync_reset;
check_mem(1364,"000011010","010000100",3,'1'); -- (0, 2, 0, 0, 1, 1, 2, 1, 0)
sync_reset;
check_mem(1365,"000011010","010000101",3,'1'); -- (0, 2, 0, 0, 1, 1, 2, 1, 2)
sync_reset;
check_mem(1366,"000011001","010000110",0,'1'); -- (0, 2, 0, 0, 1, 1, 2, 2, 1)
sync_reset;
check_mem(1367,"000010001","010001000",0,'1'); -- (0, 2, 0, 0, 1, 2, 0, 0, 1)
sync_reset;
check_mem(1368,"000010010","010001000",6,'1'); -- (0, 2, 0, 0, 1, 2, 0, 1, 0)
sync_reset;
check_mem(1369,"000010011","010001000",0,'1'); -- (0, 2, 0, 0, 1, 2, 0, 1, 1)
sync_reset;
check_mem(1370,"000010100","010001000",0,'1'); -- (0, 2, 0, 0, 1, 2, 1, 0, 0)
sync_reset;
check_mem(1371,"000010101","010001000",0,'1'); -- (0, 2, 0, 0, 1, 2, 1, 0, 1)
sync_reset;
check_mem(1372,"000010110","010001000",0,'1'); -- (0, 2, 0, 0, 1, 2, 1, 1, 0)
sync_reset;
check_mem(1373,"000010110","010001001",2,'1'); -- (0, 2, 0, 0, 1, 2, 1, 1, 2)
sync_reset;
check_mem(1374,"000010101","010001010",0,'1'); -- (0, 2, 0, 0, 1, 2, 1, 2, 1)
sync_reset;
check_mem(1375,"000010011","010001100",0,'1'); -- (0, 2, 0, 0, 1, 2, 2, 1, 1)
sync_reset;
check_mem(1376,"000000011","010010000",2,'1'); -- (0, 2, 0, 0, 2, 0, 0, 1, 1)
sync_reset;
check_mem(1377,"000000101","010010000",7,'1'); -- (0, 2, 0, 0, 2, 0, 1, 0, 1)
sync_reset;
check_mem(1378,"000000110","010010000",0,'1'); -- (0, 2, 0, 0, 2, 0, 1, 1, 0)
sync_reset;
check_mem(1379,"000001001","010010000",2,'1'); -- (0, 2, 0, 0, 2, 1, 0, 0, 1)
sync_reset;
check_mem(1380,"000001010","010010000",8,'1'); -- (0, 2, 0, 0, 2, 1, 0, 1, 0)
sync_reset;
check_mem(1381,"000001011","010010000",0,'1'); -- (0, 2, 0, 0, 2, 1, 0, 1, 1)
sync_reset;
check_mem(1382,"000001100","010010000",7,'1'); -- (0, 2, 0, 0, 2, 1, 1, 0, 0)
sync_reset;
check_mem(1383,"000001101","010010000",7,'1'); -- (0, 2, 0, 0, 2, 1, 1, 0, 1)
sync_reset;
check_mem(1384,"000001110","010010000",8,'1'); -- (0, 2, 0, 0, 2, 1, 1, 1, 0)
sync_reset;
check_mem(1385,"000001110","010010001",0,'1'); -- (0, 2, 0, 0, 2, 1, 1, 1, 2)
sync_reset;
check_mem(1386,"000001011","010010100",2,'1'); -- (0, 2, 0, 0, 2, 1, 2, 1, 1)
sync_reset;
check_mem(1387,"000100000","010000000",0,'1'); -- (0, 2, 0, 1, 0, 0, 0, 0, 0)
sync_reset;
check_mem(1388,"000100001","010000000",4,'1'); -- (0, 2, 0, 1, 0, 0, 0, 0, 1)
sync_reset;
check_mem(1389,"000100010","010000000",6,'1'); -- (0, 2, 0, 1, 0, 0, 0, 1, 0)
sync_reset;
check_mem(1390,"000100010","010000001",0,'1'); -- (0, 2, 0, 1, 0, 0, 0, 1, 2)
sync_reset;
check_mem(1391,"000100001","010000010",4,'1'); -- (0, 2, 0, 1, 0, 0, 0, 2, 1)
sync_reset;
check_mem(1392,"000100100","010000000",0,'1'); -- (0, 2, 0, 1, 0, 0, 1, 0, 0)
sync_reset;
check_mem(1393,"000100100","010000001",0,'1'); -- (0, 2, 0, 1, 0, 0, 1, 0, 2)
sync_reset;
check_mem(1394,"000100110","010000001",0,'1'); -- (0, 2, 0, 1, 0, 0, 1, 1, 2)
sync_reset;
check_mem(1395,"000100100","010000010",0,'1'); -- (0, 2, 0, 1, 0, 0, 1, 2, 0)
sync_reset;
check_mem(1396,"000100101","010000010",0,'1'); -- (0, 2, 0, 1, 0, 0, 1, 2, 1)
sync_reset;
check_mem(1397,"000100001","010000100",4,'1'); -- (0, 2, 0, 1, 0, 0, 2, 0, 1)
sync_reset;
check_mem(1398,"000100010","010000100",0,'1'); -- (0, 2, 0, 1, 0, 0, 2, 1, 0)
sync_reset;
check_mem(1399,"000100011","010000100",2,'1'); -- (0, 2, 0, 1, 0, 0, 2, 1, 1)
sync_reset;
check_mem(1400,"000101000","010000000",4,'1'); -- (0, 2, 0, 1, 0, 1, 0, 0, 0)
sync_reset;
check_mem(1401,"000101000","010000001",0,'1'); -- (0, 2, 0, 1, 0, 1, 0, 0, 2)
sync_reset;
check_mem(1402,"000101010","010000001",4,'1'); -- (0, 2, 0, 1, 0, 1, 0, 1, 2)
sync_reset;
check_mem(1403,"000101000","010000010",4,'1'); -- (0, 2, 0, 1, 0, 1, 0, 2, 0)
sync_reset;
check_mem(1404,"000101001","010000010",4,'1'); -- (0, 2, 0, 1, 0, 1, 0, 2, 1)
sync_reset;
check_mem(1405,"000101100","010000001",0,'1'); -- (0, 2, 0, 1, 0, 1, 1, 0, 2)
sync_reset;
check_mem(1406,"000101100","010000010",4,'1'); -- (0, 2, 0, 1, 0, 1, 1, 2, 0)
sync_reset;
check_mem(1407,"000101100","010000011",0,'1'); -- (0, 2, 0, 1, 0, 1, 1, 2, 2)
sync_reset;
check_mem(1408,"000101000","010000100",2,'1'); -- (0, 2, 0, 1, 0, 1, 2, 0, 0)
sync_reset;
check_mem(1409,"000101001","010000100",0,'1'); -- (0, 2, 0, 1, 0, 1, 2, 0, 1)
sync_reset;
check_mem(1410,"000101010","010000100",4,'1'); -- (0, 2, 0, 1, 0, 1, 2, 1, 0)
sync_reset;
check_mem(1411,"000101010","010000101",4,'1'); -- (0, 2, 0, 1, 0, 1, 2, 1, 2)
sync_reset;
check_mem(1412,"000101001","010000110",2,'1'); -- (0, 2, 0, 1, 0, 1, 2, 2, 1)
sync_reset;
check_mem(1413,"000100001","010001000",0,'1'); -- (0, 2, 0, 1, 0, 2, 0, 0, 1)
sync_reset;
check_mem(1414,"000100010","010001000",6,'1'); -- (0, 2, 0, 1, 0, 2, 0, 1, 0)
sync_reset;
check_mem(1415,"000100011","010001000",6,'1'); -- (0, 2, 0, 1, 0, 2, 0, 1, 1)
sync_reset;
check_mem(1416,"000100100","010001000",0,'1'); -- (0, 2, 0, 1, 0, 2, 1, 0, 0)
sync_reset;
check_mem(1417,"000100101","010001000",0,'1'); -- (0, 2, 0, 1, 0, 2, 1, 0, 1)
sync_reset;
check_mem(1418,"000100110","010001000",0,'1'); -- (0, 2, 0, 1, 0, 2, 1, 1, 0)
sync_reset;
check_mem(1419,"000100110","010001001",0,'1'); -- (0, 2, 0, 1, 0, 2, 1, 1, 2)
sync_reset;
check_mem(1420,"000100101","010001010",0,'1'); -- (0, 2, 0, 1, 0, 2, 1, 2, 1)
sync_reset;
check_mem(1421,"000100011","010001100",0,'1'); -- (0, 2, 0, 1, 0, 2, 2, 1, 1)
sync_reset;
check_mem(1422,"000110000","010000000",0,'1'); -- (0, 2, 0, 1, 1, 0, 0, 0, 0)
sync_reset;
check_mem(1423,"000110000","010000001",0,'1'); -- (0, 2, 0, 1, 1, 0, 0, 0, 2)
sync_reset;
check_mem(1424,"000110010","010000001",5,'1'); -- (0, 2, 0, 1, 1, 0, 0, 1, 2)
sync_reset;
check_mem(1425,"000110000","010000010",0,'1'); -- (0, 2, 0, 1, 1, 0, 0, 2, 0)
sync_reset;
check_mem(1426,"000110001","010000010",0,'1'); -- (0, 2, 0, 1, 1, 0, 0, 2, 1)
sync_reset;
check_mem(1427,"000110100","010000001",0,'1'); -- (0, 2, 0, 1, 1, 0, 1, 0, 2)
sync_reset;
check_mem(1428,"000110100","010000010",0,'1'); -- (0, 2, 0, 1, 1, 0, 1, 2, 0)
sync_reset;
check_mem(1429,"000110100","010000011",0,'1'); -- (0, 2, 0, 1, 1, 0, 1, 2, 2)
sync_reset;
check_mem(1430,"000110000","010000100",0,'1'); -- (0, 2, 0, 1, 1, 0, 2, 0, 0)
sync_reset;
check_mem(1431,"000110001","010000100",0,'1'); -- (0, 2, 0, 1, 1, 0, 2, 0, 1)
sync_reset;
check_mem(1432,"000110010","010000100",5,'1'); -- (0, 2, 0, 1, 1, 0, 2, 1, 0)
sync_reset;
check_mem(1433,"000110010","010000101",5,'1'); -- (0, 2, 0, 1, 1, 0, 2, 1, 2)
sync_reset;
check_mem(1434,"000110001","010000110",0,'1'); -- (0, 2, 0, 1, 1, 0, 2, 2, 1)
sync_reset;
check_mem(1435,"000110000","010001000",0,'1'); -- (0, 2, 0, 1, 1, 2, 0, 0, 0)
sync_reset;
check_mem(1436,"000110001","010001000",0,'1'); -- (0, 2, 0, 1, 1, 2, 0, 0, 1)
sync_reset;
check_mem(1437,"000110010","010001000",2,'1'); -- (0, 2, 0, 1, 1, 2, 0, 1, 0)
sync_reset;
check_mem(1438,"000110010","010001001",2,'1'); -- (0, 2, 0, 1, 1, 2, 0, 1, 2)
sync_reset;
check_mem(1439,"000110001","010001010",0,'1'); -- (0, 2, 0, 1, 1, 2, 0, 2, 1)
sync_reset;
check_mem(1440,"000110100","010001000",0,'1'); -- (0, 2, 0, 1, 1, 2, 1, 0, 0)
sync_reset;
check_mem(1441,"000110100","010001001",0,'1'); -- (0, 2, 0, 1, 1, 2, 1, 0, 2)
sync_reset;
check_mem(1442,"000110110","010001001",2,'1'); -- (0, 2, 0, 1, 1, 2, 1, 1, 2)
sync_reset;
check_mem(1443,"000110100","010001010",0,'1'); -- (0, 2, 0, 1, 1, 2, 1, 2, 0)
sync_reset;
check_mem(1444,"000110101","010001010",0,'1'); -- (0, 2, 0, 1, 1, 2, 1, 2, 1)
sync_reset;
check_mem(1445,"000110001","010001100",0,'1'); -- (0, 2, 0, 1, 1, 2, 2, 0, 1)
sync_reset;
check_mem(1446,"000110010","010001100",0,'1'); -- (0, 2, 0, 1, 1, 2, 2, 1, 0)
sync_reset;
check_mem(1447,"000110011","010001100",0,'1'); -- (0, 2, 0, 1, 1, 2, 2, 1, 1)
sync_reset;
check_mem(1448,"000100001","010010000",7,'1'); -- (0, 2, 0, 1, 2, 0, 0, 0, 1)
sync_reset;
check_mem(1449,"000100010","010010000",6,'1'); -- (0, 2, 0, 1, 2, 0, 0, 1, 0)
sync_reset;
check_mem(1450,"000100011","010010000",6,'1'); -- (0, 2, 0, 1, 2, 0, 0, 1, 1)
sync_reset;
check_mem(1451,"000100100","010010000",0,'1'); -- (0, 2, 0, 1, 2, 0, 1, 0, 0)
sync_reset;
check_mem(1452,"000100101","010010000",7,'1'); -- (0, 2, 0, 1, 2, 0, 1, 0, 1)
sync_reset;
check_mem(1453,"000100110","010010000",0,'1'); -- (0, 2, 0, 1, 2, 0, 1, 1, 0)
sync_reset;
check_mem(1454,"000100110","010010001",0,'1'); -- (0, 2, 0, 1, 2, 0, 1, 1, 2)
sync_reset;
check_mem(1455,"000100011","010010100",2,'1'); -- (0, 2, 0, 1, 2, 0, 2, 1, 1)
sync_reset;
check_mem(1456,"000101000","010010000",0,'1'); -- (0, 2, 0, 1, 2, 1, 0, 0, 0)
sync_reset;
check_mem(1457,"000101001","010010000",2,'1'); -- (0, 2, 0, 1, 2, 1, 0, 0, 1)
sync_reset;
check_mem(1458,"000101010","010010000",0,'1'); -- (0, 2, 0, 1, 2, 1, 0, 1, 0)
sync_reset;
check_mem(1459,"000101010","010010001",0,'1'); -- (0, 2, 0, 1, 2, 1, 0, 1, 2)
sync_reset;
check_mem(1460,"000101100","010010000",0,'1'); -- (0, 2, 0, 1, 2, 1, 1, 0, 0)
sync_reset;
check_mem(1461,"000101100","010010001",0,'1'); -- (0, 2, 0, 1, 2, 1, 1, 0, 2)
sync_reset;
check_mem(1462,"000101110","010010001",0,'1'); -- (0, 2, 0, 1, 2, 1, 1, 1, 2)
sync_reset;
check_mem(1463,"000101001","010010100",2,'1'); -- (0, 2, 0, 1, 2, 1, 2, 0, 1)
sync_reset;
check_mem(1464,"000101010","010010100",2,'1'); -- (0, 2, 0, 1, 2, 1, 2, 1, 0)
sync_reset;
check_mem(1465,"000101011","010010100",2,'1'); -- (0, 2, 0, 1, 2, 1, 2, 1, 1)
sync_reset;
check_mem(1466,"000100011","010011000",6,'1'); -- (0, 2, 0, 1, 2, 2, 0, 1, 1)
sync_reset;
check_mem(1467,"000100101","010011000",0,'1'); -- (0, 2, 0, 1, 2, 2, 1, 0, 1)
sync_reset;
check_mem(1468,"000100110","010011000",0,'1'); -- (0, 2, 0, 1, 2, 2, 1, 1, 0)
sync_reset;
check_mem(1469,"000000011","010100000",0,'1'); -- (0, 2, 0, 2, 0, 0, 0, 1, 1)
sync_reset;
check_mem(1470,"000000101","010100000",0,'1'); -- (0, 2, 0, 2, 0, 0, 1, 0, 1)
sync_reset;
check_mem(1471,"000000110","010100000",2,'1'); -- (0, 2, 0, 2, 0, 0, 1, 1, 0)
sync_reset;
check_mem(1472,"000001001","010100000",0,'1'); -- (0, 2, 0, 2, 0, 1, 0, 0, 1)
sync_reset;
check_mem(1473,"000001010","010100000",8,'1'); -- (0, 2, 0, 2, 0, 1, 0, 1, 0)
sync_reset;
check_mem(1474,"000001011","010100000",0,'1'); -- (0, 2, 0, 2, 0, 1, 0, 1, 1)
sync_reset;
check_mem(1475,"000001100","010100000",2,'1'); -- (0, 2, 0, 2, 0, 1, 1, 0, 0)
sync_reset;
check_mem(1476,"000001101","010100000",0,'1'); -- (0, 2, 0, 2, 0, 1, 1, 0, 1)
sync_reset;
check_mem(1477,"000001110","010100000",8,'1'); -- (0, 2, 0, 2, 0, 1, 1, 1, 0)
sync_reset;
check_mem(1478,"000001110","010100001",0,'1'); -- (0, 2, 0, 2, 0, 1, 1, 1, 2)
sync_reset;
check_mem(1479,"000001101","010100010",2,'1'); -- (0, 2, 0, 2, 0, 1, 1, 2, 1)
sync_reset;
check_mem(1480,"000001011","010100100",0,'1'); -- (0, 2, 0, 2, 0, 1, 2, 1, 1)
sync_reset;
check_mem(1481,"000010001","010100000",0,'1'); -- (0, 2, 0, 2, 1, 0, 0, 0, 1)
sync_reset;
check_mem(1482,"000010010","010100000",6,'1'); -- (0, 2, 0, 2, 1, 0, 0, 1, 0)
sync_reset;
check_mem(1483,"000010011","010100000",0,'1'); -- (0, 2, 0, 2, 1, 0, 0, 1, 1)
sync_reset;
check_mem(1484,"000010100","010100000",0,'1'); -- (0, 2, 0, 2, 1, 0, 1, 0, 0)
sync_reset;
check_mem(1485,"000010101","010100000",0,'1'); -- (0, 2, 0, 2, 1, 0, 1, 0, 1)
sync_reset;
check_mem(1486,"000010110","010100000",0,'1'); -- (0, 2, 0, 2, 1, 0, 1, 1, 0)
sync_reset;
check_mem(1487,"000010110","010100001",2,'1'); -- (0, 2, 0, 2, 1, 0, 1, 1, 2)
sync_reset;
check_mem(1488,"000010101","010100010",0,'1'); -- (0, 2, 0, 2, 1, 0, 1, 2, 1)
sync_reset;
check_mem(1489,"000010011","010100100",0,'1'); -- (0, 2, 0, 2, 1, 0, 2, 1, 1)
sync_reset;
check_mem(1490,"000011000","010100000",2,'1'); -- (0, 2, 0, 2, 1, 1, 0, 0, 0)
sync_reset;
check_mem(1491,"000011001","010100000",0,'1'); -- (0, 2, 0, 2, 1, 1, 0, 0, 1)
sync_reset;
check_mem(1492,"000011010","010100000",0,'1'); -- (0, 2, 0, 2, 1, 1, 0, 1, 0)
sync_reset;
check_mem(1493,"000011010","010100001",0,'1'); -- (0, 2, 0, 2, 1, 1, 0, 1, 2)
sync_reset;
check_mem(1494,"000011001","010100010",0,'1'); -- (0, 2, 0, 2, 1, 1, 0, 2, 1)
sync_reset;
check_mem(1495,"000011100","010100000",2,'1'); -- (0, 2, 0, 2, 1, 1, 1, 0, 0)
sync_reset;
check_mem(1496,"000011100","010100001",2,'1'); -- (0, 2, 0, 2, 1, 1, 1, 0, 2)
sync_reset;
check_mem(1497,"000011110","010100001",2,'1'); -- (0, 2, 0, 2, 1, 1, 1, 1, 2)
sync_reset;
check_mem(1498,"000011100","010100010",0,'1'); -- (0, 2, 0, 2, 1, 1, 1, 2, 0)
sync_reset;
check_mem(1499,"000011101","010100010",0,'1'); -- (0, 2, 0, 2, 1, 1, 1, 2, 1)
sync_reset;
check_mem(1500,"000011001","010100100",0,'1'); -- (0, 2, 0, 2, 1, 1, 2, 0, 1)
sync_reset;
check_mem(1501,"000011010","010100100",0,'1'); -- (0, 2, 0, 2, 1, 1, 2, 1, 0)
sync_reset;
check_mem(1502,"000011011","010100100",0,'1'); -- (0, 2, 0, 2, 1, 1, 2, 1, 1)
sync_reset;
check_mem(1503,"000010011","010101000",0,'1'); -- (0, 2, 0, 2, 1, 2, 0, 1, 1)
sync_reset;
check_mem(1504,"000010101","010101000",0,'1'); -- (0, 2, 0, 2, 1, 2, 1, 0, 1)
sync_reset;
check_mem(1505,"000010110","010101000",0,'1'); -- (0, 2, 0, 2, 1, 2, 1, 1, 0)
sync_reset;
check_mem(1506,"000001011","010110000",0,'1'); -- (0, 2, 0, 2, 2, 1, 0, 1, 1)
sync_reset;
check_mem(1507,"000001101","010110000",2,'1'); -- (0, 2, 0, 2, 2, 1, 1, 0, 1)
sync_reset;
check_mem(1508,"000001110","010110000",8,'1'); -- (0, 2, 0, 2, 2, 1, 1, 1, 0)
sync_reset;
check_mem(1509,"001000000","010000000",4,'1'); -- (0, 2, 1, 0, 0, 0, 0, 0, 0)
sync_reset;
check_mem(1510,"001000001","010000000",0,'1'); -- (0, 2, 1, 0, 0, 0, 0, 0, 1)
sync_reset;
check_mem(1511,"001000010","010000000",6,'1'); -- (0, 2, 1, 0, 0, 0, 0, 1, 0)
sync_reset;
check_mem(1512,"001000010","010000001",0,'1'); -- (0, 2, 1, 0, 0, 0, 0, 1, 2)
sync_reset;
check_mem(1513,"001000001","010000010",4,'1'); -- (0, 2, 1, 0, 0, 0, 0, 2, 1)
sync_reset;
check_mem(1514,"001000100","010000000",4,'1'); -- (0, 2, 1, 0, 0, 0, 1, 0, 0)
sync_reset;
check_mem(1515,"001000100","010000001",0,'1'); -- (0, 2, 1, 0, 0, 0, 1, 0, 2)
sync_reset;
check_mem(1516,"001000110","010000001",4,'1'); -- (0, 2, 1, 0, 0, 0, 1, 1, 2)
sync_reset;
check_mem(1517,"001000100","010000010",4,'1'); -- (0, 2, 1, 0, 0, 0, 1, 2, 0)
sync_reset;
check_mem(1518,"001000101","010000010",4,'1'); -- (0, 2, 1, 0, 0, 0, 1, 2, 1)
sync_reset;
check_mem(1519,"001000001","010000100",0,'1'); -- (0, 2, 1, 0, 0, 0, 2, 0, 1)
sync_reset;
check_mem(1520,"001000010","010000100",0,'1'); -- (0, 2, 1, 0, 0, 0, 2, 1, 0)
sync_reset;
check_mem(1521,"001000011","010000100",5,'1'); -- (0, 2, 1, 0, 0, 0, 2, 1, 1)
sync_reset;
check_mem(1522,"001001000","010000000",0,'1'); -- (0, 2, 1, 0, 0, 1, 0, 0, 0)
sync_reset;
check_mem(1523,"001001000","010000001",4,'1'); -- (0, 2, 1, 0, 0, 1, 0, 0, 2)
sync_reset;
check_mem(1524,"001001010","010000001",3,'1'); -- (0, 2, 1, 0, 0, 1, 0, 1, 2)
sync_reset;
check_mem(1525,"001001000","010000010",4,'1'); -- (0, 2, 1, 0, 0, 1, 0, 2, 0)
sync_reset;
check_mem(1526,"001001100","010000001",4,'1'); -- (0, 2, 1, 0, 0, 1, 1, 0, 2)
sync_reset;
check_mem(1527,"001001100","010000010",4,'1'); -- (0, 2, 1, 0, 0, 1, 1, 2, 0)
sync_reset;
check_mem(1528,"001001100","010000011",4,'1'); -- (0, 2, 1, 0, 0, 1, 1, 2, 2)
sync_reset;
check_mem(1529,"001001000","010000100",3,'1'); -- (0, 2, 1, 0, 0, 1, 2, 0, 0)
sync_reset;
check_mem(1530,"001001010","010000100",8,'1'); -- (0, 2, 1, 0, 0, 1, 2, 1, 0)
sync_reset;
check_mem(1531,"001001010","010000101",0,'1'); -- (0, 2, 1, 0, 0, 1, 2, 1, 2)
sync_reset;
check_mem(1532,"001000001","010001000",4,'1'); -- (0, 2, 1, 0, 0, 2, 0, 0, 1)
sync_reset;
check_mem(1533,"001000010","010001000",6,'1'); -- (0, 2, 1, 0, 0, 2, 0, 1, 0)
sync_reset;
check_mem(1534,"001000011","010001000",6,'1'); -- (0, 2, 1, 0, 0, 2, 0, 1, 1)
sync_reset;
check_mem(1535,"001000100","010001000",0,'1'); -- (0, 2, 1, 0, 0, 2, 1, 0, 0)
sync_reset;
check_mem(1536,"001000101","010001000",0,'1'); -- (0, 2, 1, 0, 0, 2, 1, 0, 1)
sync_reset;
check_mem(1537,"001000110","010001000",0,'1'); -- (0, 2, 1, 0, 0, 2, 1, 1, 0)
sync_reset;
check_mem(1538,"001000110","010001001",0,'1'); -- (0, 2, 1, 0, 0, 2, 1, 1, 2)
sync_reset;
check_mem(1539,"001000101","010001010",4,'1'); -- (0, 2, 1, 0, 0, 2, 1, 2, 1)
sync_reset;
check_mem(1540,"001000011","010001100",0,'1'); -- (0, 2, 1, 0, 0, 2, 2, 1, 1)
sync_reset;
check_mem(1541,"001010000","010000000",0,'1'); -- (0, 2, 1, 0, 1, 0, 0, 0, 0)
sync_reset;
check_mem(1542,"001010000","010000001",3,'1'); -- (0, 2, 1, 0, 1, 0, 0, 0, 2)
sync_reset;
check_mem(1543,"001010010","010000001",6,'1'); -- (0, 2, 1, 0, 1, 0, 0, 1, 2)
sync_reset;
check_mem(1544,"001010000","010000010",0,'1'); -- (0, 2, 1, 0, 1, 0, 0, 2, 0)
sync_reset;
check_mem(1545,"001010001","010000010",0,'1'); -- (0, 2, 1, 0, 1, 0, 0, 2, 1)
sync_reset;
check_mem(1546,"001010000","010000100",5,'1'); -- (0, 2, 1, 0, 1, 0, 2, 0, 0)
sync_reset;
check_mem(1547,"001010001","010000100",0,'1'); -- (0, 2, 1, 0, 1, 0, 2, 0, 1)
sync_reset;
check_mem(1548,"001010010","010000100",0,'1'); -- (0, 2, 1, 0, 1, 0, 2, 1, 0)
sync_reset;
check_mem(1549,"001010010","010000101",0,'1'); -- (0, 2, 1, 0, 1, 0, 2, 1, 2)
sync_reset;
check_mem(1550,"001010001","010000110",0,'1'); -- (0, 2, 1, 0, 1, 0, 2, 2, 1)
sync_reset;
check_mem(1551,"001011000","010000001",0,'1'); -- (0, 2, 1, 0, 1, 1, 0, 0, 2)
sync_reset;
check_mem(1552,"001011000","010000010",0,'1'); -- (0, 2, 1, 0, 1, 1, 0, 2, 0)
sync_reset;
check_mem(1553,"001011000","010000011",3,'1'); -- (0, 2, 1, 0, 1, 1, 0, 2, 2)
sync_reset;
check_mem(1554,"001011000","010000100",0,'1'); -- (0, 2, 1, 0, 1, 1, 2, 0, 0)
sync_reset;
check_mem(1555,"001011000","010000101",3,'1'); -- (0, 2, 1, 0, 1, 1, 2, 0, 2)
sync_reset;
check_mem(1556,"001011010","010000101",3,'1'); -- (0, 2, 1, 0, 1, 1, 2, 1, 2)
sync_reset;
check_mem(1557,"001011000","010000110",3,'1'); -- (0, 2, 1, 0, 1, 1, 2, 2, 0)
sync_reset;
check_mem(1558,"001010000","010001000",0,'1'); -- (0, 2, 1, 0, 1, 2, 0, 0, 0)
sync_reset;
check_mem(1559,"001010001","010001000",0,'1'); -- (0, 2, 1, 0, 1, 2, 0, 0, 1)
sync_reset;
check_mem(1560,"001010010","010001000",6,'1'); -- (0, 2, 1, 0, 1, 2, 0, 1, 0)
sync_reset;
check_mem(1561,"001010010","010001001",6,'1'); -- (0, 2, 1, 0, 1, 2, 0, 1, 2)
sync_reset;
check_mem(1562,"001010001","010001010",0,'1'); -- (0, 2, 1, 0, 1, 2, 0, 2, 1)
sync_reset;
check_mem(1563,"001010001","010001100",0,'1'); -- (0, 2, 1, 0, 1, 2, 2, 0, 1)
sync_reset;
check_mem(1564,"001010010","010001100",0,'1'); -- (0, 2, 1, 0, 1, 2, 2, 1, 0)
sync_reset;
check_mem(1565,"001010011","010001100",0,'1'); -- (0, 2, 1, 0, 1, 2, 2, 1, 1)
sync_reset;
check_mem(1566,"001000001","010010000",5,'1'); -- (0, 2, 1, 0, 2, 0, 0, 0, 1)
sync_reset;
check_mem(1567,"001000010","010010000",8,'1'); -- (0, 2, 1, 0, 2, 0, 0, 1, 0)
sync_reset;
check_mem(1568,"001000011","010010000",0,'1'); -- (0, 2, 1, 0, 2, 0, 0, 1, 1)
sync_reset;
check_mem(1569,"001000100","010010000",7,'1'); -- (0, 2, 1, 0, 2, 0, 1, 0, 0)
sync_reset;
check_mem(1570,"001000101","010010000",7,'1'); -- (0, 2, 1, 0, 2, 0, 1, 0, 1)
sync_reset;
check_mem(1571,"001000110","010010000",8,'1'); -- (0, 2, 1, 0, 2, 0, 1, 1, 0)
sync_reset;
check_mem(1572,"001000110","010010001",0,'1'); -- (0, 2, 1, 0, 2, 0, 1, 1, 2)
sync_reset;
check_mem(1573,"001000011","010010100",5,'1'); -- (0, 2, 1, 0, 2, 0, 2, 1, 1)
sync_reset;
check_mem(1574,"001001000","010010000",8,'1'); -- (0, 2, 1, 0, 2, 1, 0, 0, 0)
sync_reset;
check_mem(1575,"001001010","010010000",8,'1'); -- (0, 2, 1, 0, 2, 1, 0, 1, 0)
sync_reset;
check_mem(1576,"001001010","010010001",0,'1'); -- (0, 2, 1, 0, 2, 1, 0, 1, 2)
sync_reset;
check_mem(1577,"001001100","010010000",7,'1'); -- (0, 2, 1, 0, 2, 1, 1, 0, 0)
sync_reset;
check_mem(1578,"001001100","010010001",0,'1'); -- (0, 2, 1, 0, 2, 1, 1, 0, 2)
sync_reset;
check_mem(1579,"001001110","010010001",0,'1'); -- (0, 2, 1, 0, 2, 1, 1, 1, 2)
sync_reset;
check_mem(1580,"001001010","010010100",8,'1'); -- (0, 2, 1, 0, 2, 1, 2, 1, 0)
sync_reset;
check_mem(1581,"001000011","010011000",6,'1'); -- (0, 2, 1, 0, 2, 2, 0, 1, 1)
sync_reset;
check_mem(1582,"001000101","010011000",7,'1'); -- (0, 2, 1, 0, 2, 2, 1, 0, 1)
sync_reset;
check_mem(1583,"001000110","010011000",3,'1'); -- (0, 2, 1, 0, 2, 2, 1, 1, 0)
sync_reset;
check_mem(1584,"001100000","010000000",4,'1'); -- (0, 2, 1, 1, 0, 0, 0, 0, 0)
sync_reset;
check_mem(1585,"001100000","010000001",4,'1'); -- (0, 2, 1, 1, 0, 0, 0, 0, 2)
sync_reset;
check_mem(1586,"001100010","010000001",4,'1'); -- (0, 2, 1, 1, 0, 0, 0, 1, 2)
sync_reset;
check_mem(1587,"001100000","010000010",4,'1'); -- (0, 2, 1, 1, 0, 0, 0, 2, 0)
sync_reset;
check_mem(1588,"001100001","010000010",4,'1'); -- (0, 2, 1, 1, 0, 0, 0, 2, 1)
sync_reset;
check_mem(1589,"001100100","010000001",0,'1'); -- (0, 2, 1, 1, 0, 0, 1, 0, 2)
sync_reset;
check_mem(1590,"001100100","010000010",4,'1'); -- (0, 2, 1, 1, 0, 0, 1, 2, 0)
sync_reset;
check_mem(1591,"001100100","010000011",0,'1'); -- (0, 2, 1, 1, 0, 0, 1, 2, 2)
sync_reset;
check_mem(1592,"001100000","010000100",5,'1'); -- (0, 2, 1, 1, 0, 0, 2, 0, 0)
sync_reset;
check_mem(1593,"001100001","010000100",5,'1'); -- (0, 2, 1, 1, 0, 0, 2, 0, 1)
sync_reset;
check_mem(1594,"001100010","010000100",4,'1'); -- (0, 2, 1, 1, 0, 0, 2, 1, 0)
sync_reset;
check_mem(1595,"001100010","010000101",0,'1'); -- (0, 2, 1, 1, 0, 0, 2, 1, 2)
sync_reset;
check_mem(1596,"001100001","010000110",4,'1'); -- (0, 2, 1, 1, 0, 0, 2, 2, 1)
sync_reset;
check_mem(1597,"001101000","010000001",4,'1'); -- (0, 2, 1, 1, 0, 1, 0, 0, 2)
sync_reset;
check_mem(1598,"001101000","010000010",4,'1'); -- (0, 2, 1, 1, 0, 1, 0, 2, 0)
sync_reset;
check_mem(1599,"001101000","010000011",4,'1'); -- (0, 2, 1, 1, 0, 1, 0, 2, 2)
sync_reset;
check_mem(1600,"001101100","010000011",4,'1'); -- (0, 2, 1, 1, 0, 1, 1, 2, 2)
sync_reset;
check_mem(1601,"001101000","010000100",0,'1'); -- (0, 2, 1, 1, 0, 1, 2, 0, 0)
sync_reset;
check_mem(1602,"001101000","010000101",4,'1'); -- (0, 2, 1, 1, 0, 1, 2, 0, 2)
sync_reset;
check_mem(1603,"001101010","010000101",4,'1'); -- (0, 2, 1, 1, 0, 1, 2, 1, 2)
sync_reset;
check_mem(1604,"001101000","010000110",4,'1'); -- (0, 2, 1, 1, 0, 1, 2, 2, 0)
sync_reset;
check_mem(1605,"001100000","010001000",6,'1'); -- (0, 2, 1, 1, 0, 2, 0, 0, 0)
sync_reset;
check_mem(1606,"001100001","010001000",4,'1'); -- (0, 2, 1, 1, 0, 2, 0, 0, 1)
sync_reset;
check_mem(1607,"001100010","010001000",6,'1'); -- (0, 2, 1, 1, 0, 2, 0, 1, 0)
sync_reset;
check_mem(1608,"001100010","010001001",6,'1'); -- (0, 2, 1, 1, 0, 2, 0, 1, 2)
sync_reset;
check_mem(1609,"001100001","010001010",4,'1'); -- (0, 2, 1, 1, 0, 2, 0, 2, 1)
sync_reset;
check_mem(1610,"001100100","010001000",0,'1'); -- (0, 2, 1, 1, 0, 2, 1, 0, 0)
sync_reset;
check_mem(1611,"001100100","010001001",0,'1'); -- (0, 2, 1, 1, 0, 2, 1, 0, 2)
sync_reset;
check_mem(1612,"001100110","010001001",0,'1'); -- (0, 2, 1, 1, 0, 2, 1, 1, 2)
sync_reset;
check_mem(1613,"001100100","010001010",0,'1'); -- (0, 2, 1, 1, 0, 2, 1, 2, 0)
sync_reset;
check_mem(1614,"001100101","010001010",4,'1'); -- (0, 2, 1, 1, 0, 2, 1, 2, 1)
sync_reset;
check_mem(1615,"001100001","010001100",0,'1'); -- (0, 2, 1, 1, 0, 2, 2, 0, 1)
sync_reset;
check_mem(1616,"001100010","010001100",0,'1'); -- (0, 2, 1, 1, 0, 2, 2, 1, 0)
sync_reset;
check_mem(1617,"001100011","010001100",0,'1'); -- (0, 2, 1, 1, 0, 2, 2, 1, 1)
sync_reset;
check_mem(1618,"001110000","010000001",0,'1'); -- (0, 2, 1, 1, 1, 0, 0, 0, 2)
sync_reset;
check_mem(1619,"001110000","010000010",0,'1'); -- (0, 2, 1, 1, 1, 0, 0, 2, 0)
sync_reset;
check_mem(1620,"001110000","010000011",5,'1'); -- (0, 2, 1, 1, 1, 0, 0, 2, 2)
sync_reset;
check_mem(1621,"001110000","010000100",5,'1'); -- (0, 2, 1, 1, 1, 0, 2, 0, 0)
sync_reset;
check_mem(1622,"001110000","010000101",5,'1'); -- (0, 2, 1, 1, 1, 0, 2, 0, 2)
sync_reset;
check_mem(1623,"001110010","010000101",5,'1'); -- (0, 2, 1, 1, 1, 0, 2, 1, 2)
sync_reset;
check_mem(1624,"001110000","010000110",5,'1'); -- (0, 2, 1, 1, 1, 0, 2, 2, 0)
sync_reset;
check_mem(1625,"001110001","010000110",0,'1'); -- (0, 2, 1, 1, 1, 0, 2, 2, 1)
sync_reset;
check_mem(1626,"001110000","010001000",6,'1'); -- (0, 2, 1, 1, 1, 2, 0, 0, 0)
sync_reset;
check_mem(1627,"001110000","010001001",6,'1'); -- (0, 2, 1, 1, 1, 2, 0, 0, 2)
sync_reset;
check_mem(1628,"001110010","010001001",6,'1'); -- (0, 2, 1, 1, 1, 2, 0, 1, 2)
sync_reset;
check_mem(1629,"001110000","010001010",0,'1'); -- (0, 2, 1, 1, 1, 2, 0, 2, 0)
sync_reset;
check_mem(1630,"001110001","010001010",0,'1'); -- (0, 2, 1, 1, 1, 2, 0, 2, 1)
sync_reset;
check_mem(1631,"001110000","010001100",0,'1'); -- (0, 2, 1, 1, 1, 2, 2, 0, 0)
sync_reset;
check_mem(1632,"001110001","010001100",0,'1'); -- (0, 2, 1, 1, 1, 2, 2, 0, 1)
sync_reset;
check_mem(1633,"001110010","010001100",0,'1'); -- (0, 2, 1, 1, 1, 2, 2, 1, 0)
sync_reset;
check_mem(1634,"001110010","010001101",0,'1'); -- (0, 2, 1, 1, 1, 2, 2, 1, 2)
sync_reset;
check_mem(1635,"001110001","010001110",0,'1'); -- (0, 2, 1, 1, 1, 2, 2, 2, 1)
sync_reset;
check_mem(1636,"001100000","010010000",7,'1'); -- (0, 2, 1, 1, 2, 0, 0, 0, 0)
sync_reset;
check_mem(1637,"001100001","010010000",7,'1'); -- (0, 2, 1, 1, 2, 0, 0, 0, 1)
sync_reset;
check_mem(1638,"001100010","010010000",6,'1'); -- (0, 2, 1, 1, 2, 0, 0, 1, 0)
sync_reset;
check_mem(1639,"001100010","010010001",0,'1'); -- (0, 2, 1, 1, 2, 0, 0, 1, 2)
sync_reset;
check_mem(1640,"001100100","010010000",0,'1'); -- (0, 2, 1, 1, 2, 0, 1, 0, 0)
sync_reset;
check_mem(1641,"001100100","010010001",0,'1'); -- (0, 2, 1, 1, 2, 0, 1, 0, 2)
sync_reset;
check_mem(1642,"001100110","010010001",0,'1'); -- (0, 2, 1, 1, 2, 0, 1, 1, 2)
sync_reset;
check_mem(1643,"001100001","010010100",5,'1'); -- (0, 2, 1, 1, 2, 0, 2, 0, 1)
sync_reset;
check_mem(1644,"001100010","010010100",0,'1'); -- (0, 2, 1, 1, 2, 0, 2, 1, 0)
sync_reset;
check_mem(1645,"001100011","010010100",5,'1'); -- (0, 2, 1, 1, 2, 0, 2, 1, 1)
sync_reset;
check_mem(1646,"001101000","010010000",7,'1'); -- (0, 2, 1, 1, 2, 1, 0, 0, 0)
sync_reset;
check_mem(1647,"001101000","010010001",0,'1'); -- (0, 2, 1, 1, 2, 1, 0, 0, 2)
sync_reset;
check_mem(1648,"001101010","010010001",0,'1'); -- (0, 2, 1, 1, 2, 1, 0, 1, 2)
sync_reset;
check_mem(1649,"001101100","010010001",0,'1'); -- (0, 2, 1, 1, 2, 1, 1, 0, 2)
sync_reset;
check_mem(1650,"001101000","010010100",8,'1'); -- (0, 2, 1, 1, 2, 1, 2, 0, 0)
sync_reset;
check_mem(1651,"001101010","010010100",8,'1'); -- (0, 2, 1, 1, 2, 1, 2, 1, 0)
sync_reset;
check_mem(1652,"001101010","010010101",0,'1'); -- (0, 2, 1, 1, 2, 1, 2, 1, 2)
sync_reset;
check_mem(1653,"001100001","010011000",7,'1'); -- (0, 2, 1, 1, 2, 2, 0, 0, 1)
sync_reset;
check_mem(1654,"001100010","010011000",6,'1'); -- (0, 2, 1, 1, 2, 2, 0, 1, 0)
sync_reset;
check_mem(1655,"001100011","010011000",6,'1'); -- (0, 2, 1, 1, 2, 2, 0, 1, 1)
sync_reset;
check_mem(1656,"001100100","010011000",0,'1'); -- (0, 2, 1, 1, 2, 2, 1, 0, 0)
sync_reset;
check_mem(1657,"001100101","010011000",7,'1'); -- (0, 2, 1, 1, 2, 2, 1, 0, 1)
sync_reset;
check_mem(1658,"001100110","010011000",0,'1'); -- (0, 2, 1, 1, 2, 2, 1, 1, 0)
sync_reset;
check_mem(1659,"001100110","010011001",0,'1'); -- (0, 2, 1, 1, 2, 2, 1, 1, 2)
sync_reset;
check_mem(1660,"001100011","010011100",0,'1'); -- (0, 2, 1, 1, 2, 2, 2, 1, 1)
sync_reset;
check_mem(1661,"001000001","010100000",0,'1'); -- (0, 2, 1, 2, 0, 0, 0, 0, 1)
sync_reset;
check_mem(1662,"001000010","010100000",6,'1'); -- (0, 2, 1, 2, 0, 0, 0, 1, 0)
sync_reset;
check_mem(1663,"001000011","010100000",0,'1'); -- (0, 2, 1, 2, 0, 0, 0, 1, 1)
sync_reset;
check_mem(1664,"001000100","010100000",4,'1'); -- (0, 2, 1, 2, 0, 0, 1, 0, 0)
sync_reset;
check_mem(1665,"001000101","010100000",0,'1'); -- (0, 2, 1, 2, 0, 0, 1, 0, 1)
sync_reset;
check_mem(1666,"001000110","010100000",0,'1'); -- (0, 2, 1, 2, 0, 0, 1, 1, 0)
sync_reset;
check_mem(1667,"001000110","010100001",4,'1'); -- (0, 2, 1, 2, 0, 0, 1, 1, 2)
sync_reset;
check_mem(1668,"001000101","010100010",4,'1'); -- (0, 2, 1, 2, 0, 0, 1, 2, 1)
sync_reset;
check_mem(1669,"001000011","010100100",0,'1'); -- (0, 2, 1, 2, 0, 0, 2, 1, 1)
sync_reset;
check_mem(1670,"001001000","010100000",4,'1'); -- (0, 2, 1, 2, 0, 1, 0, 0, 0)
sync_reset;
check_mem(1671,"001001010","010100000",8,'1'); -- (0, 2, 1, 2, 0, 1, 0, 1, 0)
sync_reset;
check_mem(1672,"001001010","010100001",0,'1'); -- (0, 2, 1, 2, 0, 1, 0, 1, 2)
sync_reset;
check_mem(1673,"001001100","010100000",0,'1'); -- (0, 2, 1, 2, 0, 1, 1, 0, 0)
sync_reset;
check_mem(1674,"001001100","010100001",4,'1'); -- (0, 2, 1, 2, 0, 1, 1, 0, 2)
sync_reset;
check_mem(1675,"001001110","010100001",4,'1'); -- (0, 2, 1, 2, 0, 1, 1, 1, 2)
sync_reset;
check_mem(1676,"001001100","010100010",4,'1'); -- (0, 2, 1, 2, 0, 1, 1, 2, 0)
sync_reset;
check_mem(1677,"001001010","010100100",8,'1'); -- (0, 2, 1, 2, 0, 1, 2, 1, 0)
sync_reset;
check_mem(1678,"001000011","010101000",4,'1'); -- (0, 2, 1, 2, 0, 2, 0, 1, 1)
sync_reset;
check_mem(1679,"001000101","010101000",4,'1'); -- (0, 2, 1, 2, 0, 2, 1, 0, 1)
sync_reset;
check_mem(1680,"001000110","010101000",4,'1'); -- (0, 2, 1, 2, 0, 2, 1, 1, 0)
sync_reset;
check_mem(1681,"001010000","010100000",0,'1'); -- (0, 2, 1, 2, 1, 0, 0, 0, 0)
sync_reset;
check_mem(1682,"001010001","010100000",0,'1'); -- (0, 2, 1, 2, 1, 0, 0, 0, 1)
sync_reset;
check_mem(1683,"001010010","010100000",6,'1'); -- (0, 2, 1, 2, 1, 0, 0, 1, 0)
sync_reset;
check_mem(1684,"001010010","010100001",6,'1'); -- (0, 2, 1, 2, 1, 0, 0, 1, 2)
sync_reset;
check_mem(1685,"001010001","010100010",0,'1'); -- (0, 2, 1, 2, 1, 0, 0, 2, 1)
sync_reset;
check_mem(1686,"001010001","010100100",0,'1'); -- (0, 2, 1, 2, 1, 0, 2, 0, 1)
sync_reset;
check_mem(1687,"001010010","010100100",0,'1'); -- (0, 2, 1, 2, 1, 0, 2, 1, 0)
sync_reset;
check_mem(1688,"001010011","010100100",0,'1'); -- (0, 2, 1, 2, 1, 0, 2, 1, 1)
sync_reset;
check_mem(1689,"001011000","010100000",0,'1'); -- (0, 2, 1, 2, 1, 1, 0, 0, 0)
sync_reset;
check_mem(1690,"001011000","010100001",6,'1'); -- (0, 2, 1, 2, 1, 1, 0, 0, 2)
sync_reset;
check_mem(1691,"001011010","010100001",6,'1'); -- (0, 2, 1, 2, 1, 1, 0, 1, 2)
sync_reset;
check_mem(1692,"001011000","010100010",0,'1'); -- (0, 2, 1, 2, 1, 1, 0, 2, 0)
sync_reset;
check_mem(1693,"001011000","010100100",8,'1'); -- (0, 2, 1, 2, 1, 1, 2, 0, 0)
sync_reset;
check_mem(1694,"001011010","010100100",0,'1'); -- (0, 2, 1, 2, 1, 1, 2, 1, 0)
sync_reset;
check_mem(1695,"001011010","010100101",0,'1'); -- (0, 2, 1, 2, 1, 1, 2, 1, 2)
sync_reset;
check_mem(1696,"001010001","010101000",0,'1'); -- (0, 2, 1, 2, 1, 2, 0, 0, 1)
sync_reset;
check_mem(1697,"001010010","010101000",0,'1'); -- (0, 2, 1, 2, 1, 2, 0, 1, 0)
sync_reset;
check_mem(1698,"001010011","010101000",0,'1'); -- (0, 2, 1, 2, 1, 2, 0, 1, 1)
sync_reset;
check_mem(1699,"001010011","010101100",0,'1'); -- (0, 2, 1, 2, 1, 2, 2, 1, 1)
sync_reset;
check_mem(1700,"001000011","010110000",5,'1'); -- (0, 2, 1, 2, 2, 0, 0, 1, 1)
sync_reset;
check_mem(1701,"001000101","010110000",5,'1'); -- (0, 2, 1, 2, 2, 0, 1, 0, 1)
sync_reset;
check_mem(1702,"001000110","010110000",8,'1'); -- (0, 2, 1, 2, 2, 0, 1, 1, 0)
sync_reset;
check_mem(1703,"001001010","010110000",8,'1'); -- (0, 2, 1, 2, 2, 1, 0, 1, 0)
sync_reset;
check_mem(1704,"001001100","010110000",8,'1'); -- (0, 2, 1, 2, 2, 1, 1, 0, 0)
sync_reset;
check_mem(1705,"001001110","010110000",8,'1'); -- (0, 2, 1, 2, 2, 1, 1, 1, 0)
sync_reset;
check_mem(1706,"001001110","010110001",0,'1'); -- (0, 2, 1, 2, 2, 1, 1, 1, 2)
sync_reset;
check_mem(1707,"000000011","011000000",0,'1'); -- (0, 2, 2, 0, 0, 0, 0, 1, 1)
sync_reset;
check_mem(1708,"000000101","011000000",0,'1'); -- (0, 2, 2, 0, 0, 0, 1, 0, 1)
sync_reset;
check_mem(1709,"000000110","011000000",0,'1'); -- (0, 2, 2, 0, 0, 0, 1, 1, 0)
sync_reset;
check_mem(1710,"000001001","011000000",0,'1'); -- (0, 2, 2, 0, 0, 1, 0, 0, 1)
sync_reset;
check_mem(1711,"000001010","011000000",0,'1'); -- (0, 2, 2, 0, 0, 1, 0, 1, 0)
sync_reset;
check_mem(1712,"000001011","011000000",0,'1'); -- (0, 2, 2, 0, 0, 1, 0, 1, 1)
sync_reset;
check_mem(1713,"000001100","011000000",0,'1'); -- (0, 2, 2, 0, 0, 1, 1, 0, 0)
sync_reset;
check_mem(1714,"000001101","011000000",0,'1'); -- (0, 2, 2, 0, 0, 1, 1, 0, 1)
sync_reset;
check_mem(1715,"000001110","011000000",0,'1'); -- (0, 2, 2, 0, 0, 1, 1, 1, 0)
sync_reset;
check_mem(1716,"000001110","011000001",0,'1'); -- (0, 2, 2, 0, 0, 1, 1, 1, 2)
sync_reset;
check_mem(1717,"000001101","011000010",0,'1'); -- (0, 2, 2, 0, 0, 1, 1, 2, 1)
sync_reset;
check_mem(1718,"000001011","011000100",0,'1'); -- (0, 2, 2, 0, 0, 1, 2, 1, 1)
sync_reset;
check_mem(1719,"000010001","011000000",0,'1'); -- (0, 2, 2, 0, 1, 0, 0, 0, 1)
sync_reset;
check_mem(1720,"000010010","011000000",0,'1'); -- (0, 2, 2, 0, 1, 0, 0, 1, 0)
sync_reset;
check_mem(1721,"000010011","011000000",0,'1'); -- (0, 2, 2, 0, 1, 0, 0, 1, 1)
sync_reset;
check_mem(1722,"000010100","011000000",0,'1'); -- (0, 2, 2, 0, 1, 0, 1, 0, 0)
sync_reset;
check_mem(1723,"000010101","011000000",0,'1'); -- (0, 2, 2, 0, 1, 0, 1, 0, 1)
sync_reset;
check_mem(1724,"000010110","011000000",0,'1'); -- (0, 2, 2, 0, 1, 0, 1, 1, 0)
sync_reset;
check_mem(1725,"000010110","011000001",0,'1'); -- (0, 2, 2, 0, 1, 0, 1, 1, 2)
sync_reset;
check_mem(1726,"000010101","011000010",0,'1'); -- (0, 2, 2, 0, 1, 0, 1, 2, 1)
sync_reset;
check_mem(1727,"000010011","011000100",0,'1'); -- (0, 2, 2, 0, 1, 0, 2, 1, 1)
sync_reset;
check_mem(1728,"000011000","011000000",0,'1'); -- (0, 2, 2, 0, 1, 1, 0, 0, 0)
sync_reset;
check_mem(1729,"000011001","011000000",0,'1'); -- (0, 2, 2, 0, 1, 1, 0, 0, 1)
sync_reset;
check_mem(1730,"000011010","011000000",0,'1'); -- (0, 2, 2, 0, 1, 1, 0, 1, 0)
sync_reset;
check_mem(1731,"000011010","011000001",3,'1'); -- (0, 2, 2, 0, 1, 1, 0, 1, 2)
sync_reset;
check_mem(1732,"000011001","011000010",0,'1'); -- (0, 2, 2, 0, 1, 1, 0, 2, 1)
sync_reset;
check_mem(1733,"000011100","011000000",0,'1'); -- (0, 2, 2, 0, 1, 1, 1, 0, 0)
sync_reset;
check_mem(1734,"000011100","011000001",3,'1'); -- (0, 2, 2, 0, 1, 1, 1, 0, 2)
sync_reset;
check_mem(1735,"000011110","011000001",0,'1'); -- (0, 2, 2, 0, 1, 1, 1, 1, 2)
sync_reset;
check_mem(1736,"000011100","011000010",0,'1'); -- (0, 2, 2, 0, 1, 1, 1, 2, 0)
sync_reset;
check_mem(1737,"000011101","011000010",0,'1'); -- (0, 2, 2, 0, 1, 1, 1, 2, 1)
sync_reset;
check_mem(1738,"000011001","011000100",0,'1'); -- (0, 2, 2, 0, 1, 1, 2, 0, 1)
sync_reset;
check_mem(1739,"000011010","011000100",0,'1'); -- (0, 2, 2, 0, 1, 1, 2, 1, 0)
sync_reset;
check_mem(1740,"000011011","011000100",0,'1'); -- (0, 2, 2, 0, 1, 1, 2, 1, 1)
sync_reset;
check_mem(1741,"000010011","011001000",0,'1'); -- (0, 2, 2, 0, 1, 2, 0, 1, 1)
sync_reset;
check_mem(1742,"000010101","011001000",0,'1'); -- (0, 2, 2, 0, 1, 2, 1, 0, 1)
sync_reset;
check_mem(1743,"000010110","011001000",8,'1'); -- (0, 2, 2, 0, 1, 2, 1, 1, 0)
sync_reset;
check_mem(1744,"000001011","011010000",6,'1'); -- (0, 2, 2, 0, 2, 1, 0, 1, 1)
sync_reset;
check_mem(1745,"000001101","011010000",7,'1'); -- (0, 2, 2, 0, 2, 1, 1, 0, 1)
sync_reset;
check_mem(1746,"000001110","011010000",0,'1'); -- (0, 2, 2, 0, 2, 1, 1, 1, 0)
sync_reset;
check_mem(1747,"000100001","011000000",0,'1'); -- (0, 2, 2, 1, 0, 0, 0, 0, 1)
sync_reset;
check_mem(1748,"000100010","011000000",0,'1'); -- (0, 2, 2, 1, 0, 0, 0, 1, 0)
sync_reset;
check_mem(1749,"000100011","011000000",0,'1'); -- (0, 2, 2, 1, 0, 0, 0, 1, 1)
sync_reset;
check_mem(1750,"000100100","011000000",0,'1'); -- (0, 2, 2, 1, 0, 0, 1, 0, 0)
sync_reset;
check_mem(1751,"000100101","011000000",0,'1'); -- (0, 2, 2, 1, 0, 0, 1, 0, 1)
sync_reset;
check_mem(1752,"000100110","011000000",0,'1'); -- (0, 2, 2, 1, 0, 0, 1, 1, 0)
sync_reset;
check_mem(1753,"000100110","011000001",0,'1'); -- (0, 2, 2, 1, 0, 0, 1, 1, 2)
sync_reset;
check_mem(1754,"000100101","011000010",0,'1'); -- (0, 2, 2, 1, 0, 0, 1, 2, 1)
sync_reset;
check_mem(1755,"000100011","011000100",0,'1'); -- (0, 2, 2, 1, 0, 0, 2, 1, 1)
sync_reset;
check_mem(1756,"000101000","011000000",0,'1'); -- (0, 2, 2, 1, 0, 1, 0, 0, 0)
sync_reset;
check_mem(1757,"000101001","011000000",0,'1'); -- (0, 2, 2, 1, 0, 1, 0, 0, 1)
sync_reset;
check_mem(1758,"000101010","011000000",0,'1'); -- (0, 2, 2, 1, 0, 1, 0, 1, 0)
sync_reset;
check_mem(1759,"000101010","011000001",0,'1'); -- (0, 2, 2, 1, 0, 1, 0, 1, 2)
sync_reset;
check_mem(1760,"000101001","011000010",4,'1'); -- (0, 2, 2, 1, 0, 1, 0, 2, 1)
sync_reset;
check_mem(1761,"000101100","011000000",0,'1'); -- (0, 2, 2, 1, 0, 1, 1, 0, 0)
sync_reset;
check_mem(1762,"000101100","011000001",0,'1'); -- (0, 2, 2, 1, 0, 1, 1, 0, 2)
sync_reset;
check_mem(1763,"000101110","011000001",0,'1'); -- (0, 2, 2, 1, 0, 1, 1, 1, 2)
sync_reset;
check_mem(1764,"000101100","011000010",0,'1'); -- (0, 2, 2, 1, 0, 1, 1, 2, 0)
sync_reset;
check_mem(1765,"000101101","011000010",0,'1'); -- (0, 2, 2, 1, 0, 1, 1, 2, 1)
sync_reset;
check_mem(1766,"000101001","011000100",4,'1'); -- (0, 2, 2, 1, 0, 1, 2, 0, 1)
sync_reset;
check_mem(1767,"000101010","011000100",4,'1'); -- (0, 2, 2, 1, 0, 1, 2, 1, 0)
sync_reset;
check_mem(1768,"000101011","011000100",0,'1'); -- (0, 2, 2, 1, 0, 1, 2, 1, 1)
sync_reset;
check_mem(1769,"000100011","011001000",0,'1'); -- (0, 2, 2, 1, 0, 2, 0, 1, 1)
sync_reset;
check_mem(1770,"000100101","011001000",0,'1'); -- (0, 2, 2, 1, 0, 2, 1, 0, 1)
sync_reset;
check_mem(1771,"000100110","011001000",0,'1'); -- (0, 2, 2, 1, 0, 2, 1, 1, 0)
sync_reset;
check_mem(1772,"000110000","011000000",0,'1'); -- (0, 2, 2, 1, 1, 0, 0, 0, 0)
sync_reset;
check_mem(1773,"000110001","011000000",0,'1'); -- (0, 2, 2, 1, 1, 0, 0, 0, 1)
sync_reset;
check_mem(1774,"000110010","011000000",0,'1'); -- (0, 2, 2, 1, 1, 0, 0, 1, 0)
sync_reset;
check_mem(1775,"000110010","011000001",5,'1'); -- (0, 2, 2, 1, 1, 0, 0, 1, 2)
sync_reset;
check_mem(1776,"000110001","011000010",0,'1'); -- (0, 2, 2, 1, 1, 0, 0, 2, 1)
sync_reset;
check_mem(1777,"000110100","011000000",0,'1'); -- (0, 2, 2, 1, 1, 0, 1, 0, 0)
sync_reset;
check_mem(1778,"000110100","011000001",0,'1'); -- (0, 2, 2, 1, 1, 0, 1, 0, 2)
sync_reset;
check_mem(1779,"000110110","011000001",0,'1'); -- (0, 2, 2, 1, 1, 0, 1, 1, 2)
sync_reset;
check_mem(1780,"000110100","011000010",0,'1'); -- (0, 2, 2, 1, 1, 0, 1, 2, 0)
sync_reset;
check_mem(1781,"000110101","011000010",0,'1'); -- (0, 2, 2, 1, 1, 0, 1, 2, 1)
sync_reset;
check_mem(1782,"000110001","011000100",0,'1'); -- (0, 2, 2, 1, 1, 0, 2, 0, 1)
sync_reset;
check_mem(1783,"000110010","011000100",0,'1'); -- (0, 2, 2, 1, 1, 0, 2, 1, 0)
sync_reset;
check_mem(1784,"000110011","011000100",0,'1'); -- (0, 2, 2, 1, 1, 0, 2, 1, 1)
sync_reset;
check_mem(1785,"000110001","011001000",0,'1'); -- (0, 2, 2, 1, 1, 2, 0, 0, 1)
sync_reset;
check_mem(1786,"000110010","011001000",0,'1'); -- (0, 2, 2, 1, 1, 2, 0, 1, 0)
sync_reset;
check_mem(1787,"000110011","011001000",0,'1'); -- (0, 2, 2, 1, 1, 2, 0, 1, 1)
sync_reset;
check_mem(1788,"000110100","011001000",0,'1'); -- (0, 2, 2, 1, 1, 2, 1, 0, 0)
sync_reset;
check_mem(1789,"000110101","011001000",0,'1'); -- (0, 2, 2, 1, 1, 2, 1, 0, 1)
sync_reset;
check_mem(1790,"000110110","011001000",0,'1'); -- (0, 2, 2, 1, 1, 2, 1, 1, 0)
sync_reset;
check_mem(1791,"000110101","011001010",0,'1'); -- (0, 2, 2, 1, 1, 2, 1, 2, 1)
sync_reset;
check_mem(1792,"000110011","011001100",0,'1'); -- (0, 2, 2, 1, 1, 2, 2, 1, 1)
sync_reset;
check_mem(1793,"000100011","011010000",6,'1'); -- (0, 2, 2, 1, 2, 0, 0, 1, 1)
sync_reset;
check_mem(1794,"000100101","011010000",0,'1'); -- (0, 2, 2, 1, 2, 0, 1, 0, 1)
sync_reset;
check_mem(1795,"000100110","011010000",0,'1'); -- (0, 2, 2, 1, 2, 0, 1, 1, 0)
sync_reset;
check_mem(1796,"000101001","011010000",0,'1'); -- (0, 2, 2, 1, 2, 1, 0, 0, 1)
sync_reset;
check_mem(1797,"000101010","011010000",0,'1'); -- (0, 2, 2, 1, 2, 1, 0, 1, 0)
sync_reset;
check_mem(1798,"000101011","011010000",0,'1'); -- (0, 2, 2, 1, 2, 1, 0, 1, 1)
sync_reset;
check_mem(1799,"000101100","011010000",0,'1'); -- (0, 2, 2, 1, 2, 1, 1, 0, 0)
sync_reset;
check_mem(1800,"000101101","011010000",0,'1'); -- (0, 2, 2, 1, 2, 1, 1, 0, 1)
sync_reset;
check_mem(1801,"000101110","011010000",0,'1'); -- (0, 2, 2, 1, 2, 1, 1, 1, 0)
sync_reset;
check_mem(1802,"000101110","011010001",0,'1'); -- (0, 2, 2, 1, 2, 1, 1, 1, 2)
sync_reset;
check_mem(1803,"000001011","011100000",0,'1'); -- (0, 2, 2, 2, 0, 1, 0, 1, 1)
sync_reset;
check_mem(1804,"000001101","011100000",0,'1'); -- (0, 2, 2, 2, 0, 1, 1, 0, 1)
sync_reset;
check_mem(1805,"000001110","011100000",8,'1'); -- (0, 2, 2, 2, 0, 1, 1, 1, 0)
sync_reset;
check_mem(1806,"000010011","011100000",0,'1'); -- (0, 2, 2, 2, 1, 0, 0, 1, 1)
sync_reset;
check_mem(1807,"000010101","011100000",0,'1'); -- (0, 2, 2, 2, 1, 0, 1, 0, 1)
sync_reset;
check_mem(1808,"000010110","011100000",8,'1'); -- (0, 2, 2, 2, 1, 0, 1, 1, 0)
sync_reset;
check_mem(1809,"000011001","011100000",0,'1'); -- (0, 2, 2, 2, 1, 1, 0, 0, 1)
sync_reset;
check_mem(1810,"000011010","011100000",0,'1'); -- (0, 2, 2, 2, 1, 1, 0, 1, 0)
sync_reset;
check_mem(1811,"000011011","011100000",0,'1'); -- (0, 2, 2, 2, 1, 1, 0, 1, 1)
sync_reset;
check_mem(1812,"000011100","011100000",0,'1'); -- (0, 2, 2, 2, 1, 1, 1, 0, 0)
sync_reset;
check_mem(1813,"000011101","011100000",0,'1'); -- (0, 2, 2, 2, 1, 1, 1, 0, 1)
sync_reset;
check_mem(1814,"000011110","011100000",0,'1'); -- (0, 2, 2, 2, 1, 1, 1, 1, 0)
sync_reset;
check_mem(1815,"000011110","011100001",0,'1'); -- (0, 2, 2, 2, 1, 1, 1, 1, 2)
sync_reset;
check_mem(1816,"000011101","011100010",0,'1'); -- (0, 2, 2, 2, 1, 1, 1, 2, 1)
sync_reset;
check_mem(1817,"000011011","011100100",0,'1'); -- (0, 2, 2, 2, 1, 1, 2, 1, 1)
sync_reset;
check_mem(1818,"100000000","000000000",4,'1'); -- (1, 0, 0, 0, 0, 0, 0, 0, 0)
sync_reset;
check_mem(1819,"100000000","000000001",2,'1'); -- (1, 0, 0, 0, 0, 0, 0, 0, 2)
sync_reset;
check_mem(1820,"100000010","000000001",1,'1'); -- (1, 0, 0, 0, 0, 0, 0, 1, 2)
sync_reset;
check_mem(1821,"100000000","000000010",2,'1'); -- (1, 0, 0, 0, 0, 0, 0, 2, 0)
sync_reset;
check_mem(1822,"100000001","000000010",4,'1'); -- (1, 0, 0, 0, 0, 0, 0, 2, 1)
sync_reset;
check_mem(1823,"100000100","000000001",1,'1'); -- (1, 0, 0, 0, 0, 0, 1, 0, 2)
sync_reset;
check_mem(1824,"100000100","000000010",1,'1'); -- (1, 0, 0, 0, 0, 0, 1, 2, 0)
sync_reset;
check_mem(1825,"100000100","000000011",1,'1'); -- (1, 0, 0, 0, 0, 0, 1, 2, 2)
sync_reset;
check_mem(1826,"100000000","000000100",1,'1'); -- (1, 0, 0, 0, 0, 0, 2, 0, 0)
sync_reset;
check_mem(1827,"100000001","000000100",1,'1'); -- (1, 0, 0, 0, 0, 0, 2, 0, 1)
sync_reset;
check_mem(1828,"100000010","000000100",1,'1'); -- (1, 0, 0, 0, 0, 0, 2, 1, 0)
sync_reset;
check_mem(1829,"100000010","000000101",1,'1'); -- (1, 0, 0, 0, 0, 0, 2, 1, 2)
sync_reset;
check_mem(1830,"100000001","000000110",1,'1'); -- (1, 0, 0, 0, 0, 0, 2, 2, 1)
sync_reset;
check_mem(1831,"100001000","000000001",3,'1'); -- (1, 0, 0, 0, 0, 1, 0, 0, 2)
sync_reset;
check_mem(1832,"100001000","000000010",4,'1'); -- (1, 0, 0, 0, 0, 1, 0, 2, 0)
sync_reset;
check_mem(1833,"100001000","000000011",6,'1'); -- (1, 0, 0, 0, 0, 1, 0, 2, 2)
sync_reset;
check_mem(1834,"100001100","000000011",1,'1'); -- (1, 0, 0, 0, 0, 1, 1, 2, 2)
sync_reset;
check_mem(1835,"100001000","000000100",8,'1'); -- (1, 0, 0, 0, 0, 1, 2, 0, 0)
sync_reset;
check_mem(1836,"100001000","000000101",7,'1'); -- (1, 0, 0, 0, 0, 1, 2, 0, 2)
sync_reset;
check_mem(1837,"100001010","000000101",1,'1'); -- (1, 0, 0, 0, 0, 1, 2, 1, 2)
sync_reset;
check_mem(1838,"100001000","000000110",8,'1'); -- (1, 0, 0, 0, 0, 1, 2, 2, 0)
sync_reset;
check_mem(1839,"100001001","000000110",1,'1'); -- (1, 0, 0, 0, 0, 1, 2, 2, 1)
sync_reset;
check_mem(1840,"100000000","000001000",2,'1'); -- (1, 0, 0, 0, 0, 2, 0, 0, 0)
sync_reset;
check_mem(1841,"100000001","000001000",4,'1'); -- (1, 0, 0, 0, 0, 2, 0, 0, 1)
sync_reset;
check_mem(1842,"100000010","000001000",4,'1'); -- (1, 0, 0, 0, 0, 2, 0, 1, 0)
sync_reset;
check_mem(1843,"100000010","000001001",2,'1'); -- (1, 0, 0, 0, 0, 2, 0, 1, 2)
sync_reset;
check_mem(1844,"100000001","000001010",1,'1'); -- (1, 0, 0, 0, 0, 2, 0, 2, 1)
sync_reset;
check_mem(1845,"100000100","000001000",1,'1'); -- (1, 0, 0, 0, 0, 2, 1, 0, 0)
sync_reset;
check_mem(1846,"100000100","000001001",2,'1'); -- (1, 0, 0, 0, 0, 2, 1, 0, 2)
sync_reset;
check_mem(1847,"100000110","000001001",2,'1'); -- (1, 0, 0, 0, 0, 2, 1, 1, 2)
sync_reset;
check_mem(1848,"100000100","000001010",1,'1'); -- (1, 0, 0, 0, 0, 2, 1, 2, 0)
sync_reset;
check_mem(1849,"100000101","000001010",1,'1'); -- (1, 0, 0, 0, 0, 2, 1, 2, 1)
sync_reset;
check_mem(1850,"100000001","000001100",1,'1'); -- (1, 0, 0, 0, 0, 2, 2, 0, 1)
sync_reset;
check_mem(1851,"100000010","000001100",1,'1'); -- (1, 0, 0, 0, 0, 2, 2, 1, 0)
sync_reset;
check_mem(1852,"100000011","000001100",4,'1'); -- (1, 0, 0, 0, 0, 2, 2, 1, 1)
sync_reset;
check_mem(1853,"100010000","000000001",2,'1'); -- (1, 0, 0, 0, 1, 0, 0, 0, 2)
sync_reset;
check_mem(1854,"100010000","000000010",1,'1'); -- (1, 0, 0, 0, 1, 0, 0, 2, 0)
sync_reset;
check_mem(1855,"100010000","000000011",6,'1'); -- (1, 0, 0, 0, 1, 0, 0, 2, 2)
sync_reset;
check_mem(1856,"100010100","000000011",1,'1'); -- (1, 0, 0, 0, 1, 0, 1, 2, 2)
sync_reset;
check_mem(1857,"100010000","000000100",8,'1'); -- (1, 0, 0, 0, 1, 0, 2, 0, 0)
sync_reset;
check_mem(1858,"100010000","000000101",7,'1'); -- (1, 0, 0, 0, 1, 0, 2, 0, 2)
sync_reset;
check_mem(1859,"100010010","000000101",1,'1'); -- (1, 0, 0, 0, 1, 0, 2, 1, 2)
sync_reset;
check_mem(1860,"100010000","000000110",8,'1'); -- (1, 0, 0, 0, 1, 0, 2, 2, 0)
sync_reset;
check_mem(1861,"100011000","000000011",6,'1'); -- (1, 0, 0, 0, 1, 1, 0, 2, 2)
sync_reset;
check_mem(1862,"100011000","000000101",7,'1'); -- (1, 0, 0, 0, 1, 1, 2, 0, 2)
sync_reset;
check_mem(1863,"100011000","000000110",8,'1'); -- (1, 0, 0, 0, 1, 1, 2, 2, 0)
sync_reset;
check_mem(1864,"100010000","000001000",1,'1'); -- (1, 0, 0, 0, 1, 2, 0, 0, 0)
sync_reset;
check_mem(1865,"100010000","000001001",2,'1'); -- (1, 0, 0, 0, 1, 2, 0, 0, 2)
sync_reset;
check_mem(1866,"100010010","000001001",2,'1'); -- (1, 0, 0, 0, 1, 2, 0, 1, 2)
sync_reset;
check_mem(1867,"100010000","000001010",1,'1'); -- (1, 0, 0, 0, 1, 2, 0, 2, 0)
sync_reset;
check_mem(1868,"100010100","000001001",2,'1'); -- (1, 0, 0, 0, 1, 2, 1, 0, 2)
sync_reset;
check_mem(1869,"100010100","000001010",1,'1'); -- (1, 0, 0, 0, 1, 2, 1, 2, 0)
sync_reset;
check_mem(1870,"100010100","000001011",2,'1'); -- (1, 0, 0, 0, 1, 2, 1, 2, 2)
sync_reset;
check_mem(1871,"100010000","000001100",1,'1'); -- (1, 0, 0, 0, 1, 2, 2, 0, 0)
sync_reset;
check_mem(1872,"100010010","000001100",1,'1'); -- (1, 0, 0, 0, 1, 2, 2, 1, 0)
sync_reset;
check_mem(1873,"100010010","000001101",1,'1'); -- (1, 0, 0, 0, 1, 2, 2, 1, 2)
sync_reset;
check_mem(1874,"100000000","000010000",1,'1'); -- (1, 0, 0, 0, 2, 0, 0, 0, 0)
sync_reset;
check_mem(1875,"100000001","000010000",1,'1'); -- (1, 0, 0, 0, 2, 0, 0, 0, 1)
sync_reset;
check_mem(1876,"100000010","000010000",3,'1'); -- (1, 0, 0, 0, 2, 0, 0, 1, 0)
sync_reset;
check_mem(1877,"100000010","000010001",2,'1'); -- (1, 0, 0, 0, 2, 0, 0, 1, 2)
sync_reset;
check_mem(1878,"100000001","000010010",1,'1'); -- (1, 0, 0, 0, 2, 0, 0, 2, 1)
sync_reset;
check_mem(1879,"100000100","000010000",3,'1'); -- (1, 0, 0, 0, 2, 0, 1, 0, 0)
sync_reset;
check_mem(1880,"100000100","000010001",1,'1'); -- (1, 0, 0, 0, 2, 0, 1, 0, 2)
sync_reset;
check_mem(1881,"100000110","000010001",3,'1'); -- (1, 0, 0, 0, 2, 0, 1, 1, 2)
sync_reset;
check_mem(1882,"100000100","000010010",1,'1'); -- (1, 0, 0, 0, 2, 0, 1, 2, 0)
sync_reset;
check_mem(1883,"100000101","000010010",1,'1'); -- (1, 0, 0, 0, 2, 0, 1, 2, 1)
sync_reset;
check_mem(1884,"100000001","000010100",2,'1'); -- (1, 0, 0, 0, 2, 0, 2, 0, 1)
sync_reset;
check_mem(1885,"100000010","000010100",2,'1'); -- (1, 0, 0, 0, 2, 0, 2, 1, 0)
sync_reset;
check_mem(1886,"100000011","000010100",2,'1'); -- (1, 0, 0, 0, 2, 0, 2, 1, 1)
sync_reset;
check_mem(1887,"100001000","000010000",1,'1'); -- (1, 0, 0, 0, 2, 1, 0, 0, 0)
sync_reset;
check_mem(1888,"100001000","000010001",1,'1'); -- (1, 0, 0, 0, 2, 1, 0, 0, 2)
sync_reset;
check_mem(1889,"100001010","000010001",1,'1'); -- (1, 0, 0, 0, 2, 1, 0, 1, 2)
sync_reset;
check_mem(1890,"100001000","000010010",1,'1'); -- (1, 0, 0, 0, 2, 1, 0, 2, 0)
sync_reset;
check_mem(1891,"100001001","000010010",1,'1'); -- (1, 0, 0, 0, 2, 1, 0, 2, 1)
sync_reset;
check_mem(1892,"100001100","000010001",3,'1'); -- (1, 0, 0, 0, 2, 1, 1, 0, 2)
sync_reset;
check_mem(1893,"100001100","000010010",1,'1'); -- (1, 0, 0, 0, 2, 1, 1, 2, 0)
sync_reset;
check_mem(1894,"100001100","000010011",1,'1'); -- (1, 0, 0, 0, 2, 1, 1, 2, 2)
sync_reset;
check_mem(1895,"100001000","000010100",2,'1'); -- (1, 0, 0, 0, 2, 1, 2, 0, 0)
sync_reset;
check_mem(1896,"100001001","000010100",2,'1'); -- (1, 0, 0, 0, 2, 1, 2, 0, 1)
sync_reset;
check_mem(1897,"100001010","000010100",2,'1'); -- (1, 0, 0, 0, 2, 1, 2, 1, 0)
sync_reset;
check_mem(1898,"100001010","000010101",2,'1'); -- (1, 0, 0, 0, 2, 1, 2, 1, 2)
sync_reset;
check_mem(1899,"100001001","000010110",2,'1'); -- (1, 0, 0, 0, 2, 1, 2, 2, 1)
sync_reset;
check_mem(1900,"100000001","000011000",3,'1'); -- (1, 0, 0, 0, 2, 2, 0, 0, 1)
sync_reset;
check_mem(1901,"100000010","000011000",3,'1'); -- (1, 0, 0, 0, 2, 2, 0, 1, 0)
sync_reset;
check_mem(1902,"100000011","000011000",3,'1'); -- (1, 0, 0, 0, 2, 2, 0, 1, 1)
sync_reset;
check_mem(1903,"100000100","000011000",3,'1'); -- (1, 0, 0, 0, 2, 2, 1, 0, 0)
sync_reset;
check_mem(1904,"100000101","000011000",3,'1'); -- (1, 0, 0, 0, 2, 2, 1, 0, 1)
sync_reset;
check_mem(1905,"100000110","000011000",3,'1'); -- (1, 0, 0, 0, 2, 2, 1, 1, 0)
sync_reset;
check_mem(1906,"100000110","000011001",3,'1'); -- (1, 0, 0, 0, 2, 2, 1, 1, 2)
sync_reset;
check_mem(1907,"100000101","000011010",3,'1'); -- (1, 0, 0, 0, 2, 2, 1, 2, 1)
sync_reset;
check_mem(1908,"100000011","000011100",1,'1'); -- (1, 0, 0, 0, 2, 2, 2, 1, 1)
sync_reset;
check_mem(1909,"100100000","000000001",6,'1'); -- (1, 0, 0, 1, 0, 0, 0, 0, 2)
sync_reset;
check_mem(1910,"100100000","000000010",6,'1'); -- (1, 0, 0, 1, 0, 0, 0, 2, 0)
sync_reset;
check_mem(1911,"100100000","000000011",6,'1'); -- (1, 0, 0, 1, 0, 0, 0, 2, 2)
sync_reset;
check_mem(1912,"100100000","000000100",7,'1'); -- (1, 0, 0, 1, 0, 0, 2, 0, 0)
sync_reset;
check_mem(1913,"100100000","000000101",1,'1'); -- (1, 0, 0, 1, 0, 0, 2, 0, 2)
sync_reset;
check_mem(1914,"100100010","000000101",2,'1'); -- (1, 0, 0, 1, 0, 0, 2, 1, 2)
sync_reset;
check_mem(1915,"100100000","000000110",1,'1'); -- (1, 0, 0, 1, 0, 0, 2, 2, 0)
sync_reset;
check_mem(1916,"100100001","000000110",4,'1'); -- (1, 0, 0, 1, 0, 0, 2, 2, 1)
sync_reset;
check_mem(1917,"100101000","000000011",6,'1'); -- (1, 0, 0, 1, 0, 1, 0, 2, 2)
sync_reset;
check_mem(1918,"100101000","000000101",4,'1'); -- (1, 0, 0, 1, 0, 1, 2, 0, 2)
sync_reset;
check_mem(1919,"100101000","000000110",4,'1'); -- (1, 0, 0, 1, 0, 1, 2, 2, 0)
sync_reset;
check_mem(1920,"100100000","000001000",6,'1'); -- (1, 0, 0, 1, 0, 2, 0, 0, 0)
sync_reset;
check_mem(1921,"100100000","000001001",2,'1'); -- (1, 0, 0, 1, 0, 2, 0, 0, 2)
sync_reset;
check_mem(1922,"100100010","000001001",2,'1'); -- (1, 0, 0, 1, 0, 2, 0, 1, 2)
sync_reset;
check_mem(1923,"100100000","000001010",1,'1'); -- (1, 0, 0, 1, 0, 2, 0, 2, 0)
sync_reset;
check_mem(1924,"100100001","000001010",1,'1'); -- (1, 0, 0, 1, 0, 2, 0, 2, 1)
sync_reset;
check_mem(1925,"100100000","000001100",2,'1'); -- (1, 0, 0, 1, 0, 2, 2, 0, 0)
sync_reset;
check_mem(1926,"100100001","000001100",4,'1'); -- (1, 0, 0, 1, 0, 2, 2, 0, 1)
sync_reset;
check_mem(1927,"100100010","000001100",2,'1'); -- (1, 0, 0, 1, 0, 2, 2, 1, 0)
sync_reset;
check_mem(1928,"100100010","000001101",2,'1'); -- (1, 0, 0, 1, 0, 2, 2, 1, 2)
sync_reset;
check_mem(1929,"100100001","000001110",1,'1'); -- (1, 0, 0, 1, 0, 2, 2, 2, 1)
sync_reset;
check_mem(1930,"100110000","000000011",6,'1'); -- (1, 0, 0, 1, 1, 0, 0, 2, 2)
sync_reset;
check_mem(1931,"100110000","000000101",5,'1'); -- (1, 0, 0, 1, 1, 0, 2, 0, 2)
sync_reset;
check_mem(1932,"100110000","000000110",8,'1'); -- (1, 0, 0, 1, 1, 0, 2, 2, 0)
sync_reset;
check_mem(1933,"100110000","000001001",2,'1'); -- (1, 0, 0, 1, 1, 2, 0, 0, 2)
sync_reset;
check_mem(1934,"100110000","000001010",1,'1'); -- (1, 0, 0, 1, 1, 2, 0, 2, 0)
sync_reset;
check_mem(1935,"100110000","000001011",6,'1'); -- (1, 0, 0, 1, 1, 2, 0, 2, 2)
sync_reset;
check_mem(1936,"100110000","000001100",8,'1'); -- (1, 0, 0, 1, 1, 2, 2, 0, 0)
sync_reset;
check_mem(1937,"100110000","000001101",1,'1'); -- (1, 0, 0, 1, 1, 2, 2, 0, 2)
sync_reset;
check_mem(1938,"100110010","000001101",2,'1'); -- (1, 0, 0, 1, 1, 2, 2, 1, 2)
sync_reset;
check_mem(1939,"100110000","000001110",8,'1'); -- (1, 0, 0, 1, 1, 2, 2, 2, 0)
sync_reset;
check_mem(1940,"100100000","000010000",6,'1'); -- (1, 0, 0, 1, 2, 0, 0, 0, 0)
sync_reset;
check_mem(1941,"100100000","000010001",1,'1'); -- (1, 0, 0, 1, 2, 0, 0, 0, 2)
sync_reset;
check_mem(1942,"100100010","000010001",6,'1'); -- (1, 0, 0, 1, 2, 0, 0, 1, 2)
sync_reset;
check_mem(1943,"100100000","000010010",1,'1'); -- (1, 0, 0, 1, 2, 0, 0, 2, 0)
sync_reset;
check_mem(1944,"100100001","000010010",1,'1'); -- (1, 0, 0, 1, 2, 0, 0, 2, 1)
sync_reset;
check_mem(1945,"100100000","000010100",2,'1'); -- (1, 0, 0, 1, 2, 0, 2, 0, 0)
sync_reset;
check_mem(1946,"100100001","000010100",1,'1'); -- (1, 0, 0, 1, 2, 0, 2, 0, 1)
sync_reset;
check_mem(1947,"100100010","000010100",2,'1'); -- (1, 0, 0, 1, 2, 0, 2, 1, 0)
sync_reset;
check_mem(1948,"100100010","000010101",2,'1'); -- (1, 0, 0, 1, 2, 0, 2, 1, 2)
sync_reset;
check_mem(1949,"100100001","000010110",1,'1'); -- (1, 0, 0, 1, 2, 0, 2, 2, 1)
sync_reset;
check_mem(1950,"100101000","000010001",6,'1'); -- (1, 0, 0, 1, 2, 1, 0, 0, 2)
sync_reset;
check_mem(1951,"100101000","000010010",1,'1'); -- (1, 0, 0, 1, 2, 1, 0, 2, 0)
sync_reset;
check_mem(1952,"100101000","000010011",6,'1'); -- (1, 0, 0, 1, 2, 1, 0, 2, 2)
sync_reset;
check_mem(1953,"100101000","000010100",1,'1'); -- (1, 0, 0, 1, 2, 1, 2, 0, 0)
sync_reset;
check_mem(1954,"100101000","000010101",1,'1'); -- (1, 0, 0, 1, 2, 1, 2, 0, 2)
sync_reset;
check_mem(1955,"100101010","000010101",2,'1'); -- (1, 0, 0, 1, 2, 1, 2, 1, 2)
sync_reset;
check_mem(1956,"100101000","000010110",1,'1'); -- (1, 0, 0, 1, 2, 1, 2, 2, 0)
sync_reset;
check_mem(1957,"100101001","000010110",1,'1'); -- (1, 0, 0, 1, 2, 1, 2, 2, 1)
sync_reset;
check_mem(1958,"100100000","000011000",1,'1'); -- (1, 0, 0, 1, 2, 2, 0, 0, 0)
sync_reset;
check_mem(1959,"100100001","000011000",6,'1'); -- (1, 0, 0, 1, 2, 2, 0, 0, 1)
sync_reset;
check_mem(1960,"100100010","000011000",6,'1'); -- (1, 0, 0, 1, 2, 2, 0, 1, 0)
sync_reset;
check_mem(1961,"100100010","000011001",2,'1'); -- (1, 0, 0, 1, 2, 2, 0, 1, 2)
sync_reset;
check_mem(1962,"100100001","000011010",1,'1'); -- (1, 0, 0, 1, 2, 2, 0, 2, 1)
sync_reset;
check_mem(1963,"100100001","000011100",2,'1'); -- (1, 0, 0, 1, 2, 2, 2, 0, 1)
sync_reset;
check_mem(1964,"100100010","000011100",2,'1'); -- (1, 0, 0, 1, 2, 2, 2, 1, 0)
sync_reset;
check_mem(1965,"100100011","000011100",2,'1'); -- (1, 0, 0, 1, 2, 2, 2, 1, 1)
sync_reset;
check_mem(1966,"100000000","000100000",1,'1'); -- (1, 0, 0, 2, 0, 0, 0, 0, 0)
sync_reset;
check_mem(1967,"100000001","000100000",4,'1'); -- (1, 0, 0, 2, 0, 0, 0, 0, 1)
sync_reset;
check_mem(1968,"100000010","000100000",4,'1'); -- (1, 0, 0, 2, 0, 0, 0, 1, 0)
sync_reset;
check_mem(1969,"100000010","000100001",1,'1'); -- (1, 0, 0, 2, 0, 0, 0, 1, 2)
sync_reset;
check_mem(1970,"100000001","000100010",1,'1'); -- (1, 0, 0, 2, 0, 0, 0, 2, 1)
sync_reset;
check_mem(1971,"100000100","000100000",4,'1'); -- (1, 0, 0, 2, 0, 0, 1, 0, 0)
sync_reset;
check_mem(1972,"100000100","000100001",2,'1'); -- (1, 0, 0, 2, 0, 0, 1, 0, 2)
sync_reset;
check_mem(1973,"100000110","000100001",5,'1'); -- (1, 0, 0, 2, 0, 0, 1, 1, 2)
sync_reset;
check_mem(1974,"100000100","000100010",2,'1'); -- (1, 0, 0, 2, 0, 0, 1, 2, 0)
sync_reset;
check_mem(1975,"100000101","000100010",4,'1'); -- (1, 0, 0, 2, 0, 0, 1, 2, 1)
sync_reset;
check_mem(1976,"100000001","000100100",1,'1'); -- (1, 0, 0, 2, 0, 0, 2, 0, 1)
sync_reset;
check_mem(1977,"100000010","000100100",1,'1'); -- (1, 0, 0, 2, 0, 0, 2, 1, 0)
sync_reset;
check_mem(1978,"100000011","000100100",4,'1'); -- (1, 0, 0, 2, 0, 0, 2, 1, 1)
sync_reset;
check_mem(1979,"100001000","000100000",2,'1'); -- (1, 0, 0, 2, 0, 1, 0, 0, 0)
sync_reset;
check_mem(1980,"100001000","000100001",1,'1'); -- (1, 0, 0, 2, 0, 1, 0, 0, 2)
sync_reset;
check_mem(1981,"100001010","000100001",1,'1'); -- (1, 0, 0, 2, 0, 1, 0, 1, 2)
sync_reset;
check_mem(1982,"100001000","000100010",2,'1'); -- (1, 0, 0, 2, 0, 1, 0, 2, 0)
sync_reset;
check_mem(1983,"100001001","000100010",1,'1'); -- (1, 0, 0, 2, 0, 1, 0, 2, 1)
sync_reset;
check_mem(1984,"100001100","000100001",1,'1'); -- (1, 0, 0, 2, 0, 1, 1, 0, 2)
sync_reset;
check_mem(1985,"100001100","000100010",2,'1'); -- (1, 0, 0, 2, 0, 1, 1, 2, 0)
sync_reset;
check_mem(1986,"100001100","000100011",2,'1'); -- (1, 0, 0, 2, 0, 1, 1, 2, 2)
sync_reset;
check_mem(1987,"100001000","000100100",1,'1'); -- (1, 0, 0, 2, 0, 1, 2, 0, 0)
sync_reset;
check_mem(1988,"100001001","000100100",1,'1'); -- (1, 0, 0, 2, 0, 1, 2, 0, 1)
sync_reset;
check_mem(1989,"100001010","000100100",1,'1'); -- (1, 0, 0, 2, 0, 1, 2, 1, 0)
sync_reset;
check_mem(1990,"100001010","000100101",1,'1'); -- (1, 0, 0, 2, 0, 1, 2, 1, 2)
sync_reset;
check_mem(1991,"100001001","000100110",1,'1'); -- (1, 0, 0, 2, 0, 1, 2, 2, 1)
sync_reset;
check_mem(1992,"100000001","000101000",4,'1'); -- (1, 0, 0, 2, 0, 2, 0, 0, 1)
sync_reset;
check_mem(1993,"100000010","000101000",4,'1'); -- (1, 0, 0, 2, 0, 2, 0, 1, 0)
sync_reset;
check_mem(1994,"100000011","000101000",4,'1'); -- (1, 0, 0, 2, 0, 2, 0, 1, 1)
sync_reset;
check_mem(1995,"100000100","000101000",4,'1'); -- (1, 0, 0, 2, 0, 2, 1, 0, 0)
sync_reset;
check_mem(1996,"100000101","000101000",4,'1'); -- (1, 0, 0, 2, 0, 2, 1, 0, 1)
sync_reset;
check_mem(1997,"100000110","000101000",4,'1'); -- (1, 0, 0, 2, 0, 2, 1, 1, 0)
sync_reset;
check_mem(1998,"100000110","000101001",1,'1'); -- (1, 0, 0, 2, 0, 2, 1, 1, 2)
sync_reset;
check_mem(1999,"100000101","000101010",4,'1'); -- (1, 0, 0, 2, 0, 2, 1, 2, 1)
sync_reset;
check_mem(2000,"100000011","000101100",4,'1'); -- (1, 0, 0, 2, 0, 2, 2, 1, 1)
sync_reset;
check_mem(2001,"100010000","000100000",1,'1'); -- (1, 0, 0, 2, 1, 0, 0, 0, 0)
sync_reset;
check_mem(2002,"100010000","000100001",1,'1'); -- (1, 0, 0, 2, 1, 0, 0, 0, 2)
sync_reset;
check_mem(2003,"100010010","000100001",1,'1'); -- (1, 0, 0, 2, 1, 0, 0, 1, 2)
sync_reset;
check_mem(2004,"100010000","000100010",1,'1'); -- (1, 0, 0, 2, 1, 0, 0, 2, 0)
sync_reset;
check_mem(2005,"100010100","000100001",2,'1'); -- (1, 0, 0, 2, 1, 0, 1, 0, 2)
sync_reset;
check_mem(2006,"100010100","000100010",1,'1'); -- (1, 0, 0, 2, 1, 0, 1, 2, 0)
sync_reset;
check_mem(2007,"100010100","000100011",2,'1'); -- (1, 0, 0, 2, 1, 0, 1, 2, 2)
sync_reset;
check_mem(2008,"100010000","000100100",1,'1'); -- (1, 0, 0, 2, 1, 0, 2, 0, 0)
sync_reset;
check_mem(2009,"100010010","000100100",1,'1'); -- (1, 0, 0, 2, 1, 0, 2, 1, 0)
sync_reset;
check_mem(2010,"100010010","000100101",1,'1'); -- (1, 0, 0, 2, 1, 0, 2, 1, 2)
sync_reset;
check_mem(2011,"100011000","000100001",1,'1'); -- (1, 0, 0, 2, 1, 1, 0, 0, 2)
sync_reset;
check_mem(2012,"100011000","000100010",8,'1'); -- (1, 0, 0, 2, 1, 1, 0, 2, 0)
sync_reset;
check_mem(2013,"100011000","000100011",6,'1'); -- (1, 0, 0, 2, 1, 1, 0, 2, 2)
sync_reset;
check_mem(2014,"100011100","000100011",2,'1'); -- (1, 0, 0, 2, 1, 1, 1, 2, 2)
sync_reset;
check_mem(2015,"100011000","000100100",8,'1'); -- (1, 0, 0, 2, 1, 1, 2, 0, 0)
sync_reset;
check_mem(2016,"100011000","000100101",7,'1'); -- (1, 0, 0, 2, 1, 1, 2, 0, 2)
sync_reset;
check_mem(2017,"100011010","000100101",1,'1'); -- (1, 0, 0, 2, 1, 1, 2, 1, 2)
sync_reset;
check_mem(2018,"100011000","000100110",8,'1'); -- (1, 0, 0, 2, 1, 1, 2, 2, 0)
sync_reset;
check_mem(2019,"100010000","000101000",1,'1'); -- (1, 0, 0, 2, 1, 2, 0, 0, 0)
sync_reset;
check_mem(2020,"100010010","000101000",1,'1'); -- (1, 0, 0, 2, 1, 2, 0, 1, 0)
sync_reset;
check_mem(2021,"100010010","000101001",1,'1'); -- (1, 0, 0, 2, 1, 2, 0, 1, 2)
sync_reset;
check_mem(2022,"100010100","000101000",1,'1'); -- (1, 0, 0, 2, 1, 2, 1, 0, 0)
sync_reset;
check_mem(2023,"100010100","000101001",2,'1'); -- (1, 0, 0, 2, 1, 2, 1, 0, 2)
sync_reset;
check_mem(2024,"100010110","000101001",2,'1'); -- (1, 0, 0, 2, 1, 2, 1, 1, 2)
sync_reset;
check_mem(2025,"100010100","000101010",1,'1'); -- (1, 0, 0, 2, 1, 2, 1, 2, 0)
sync_reset;
check_mem(2026,"100010010","000101100",1,'1'); -- (1, 0, 0, 2, 1, 2, 2, 1, 0)
sync_reset;
check_mem(2027,"100000001","000110000",5,'1'); -- (1, 0, 0, 2, 2, 0, 0, 0, 1)
sync_reset;
check_mem(2028,"100000010","000110000",5,'1'); -- (1, 0, 0, 2, 2, 0, 0, 1, 0)
sync_reset;
check_mem(2029,"100000011","000110000",5,'1'); -- (1, 0, 0, 2, 2, 0, 0, 1, 1)
sync_reset;
check_mem(2030,"100000100","000110000",5,'1'); -- (1, 0, 0, 2, 2, 0, 1, 0, 0)
sync_reset;
check_mem(2031,"100000101","000110000",5,'1'); -- (1, 0, 0, 2, 2, 0, 1, 0, 1)
sync_reset;
check_mem(2032,"100000110","000110000",5,'1'); -- (1, 0, 0, 2, 2, 0, 1, 1, 0)
sync_reset;
check_mem(2033,"100000110","000110001",5,'1'); -- (1, 0, 0, 2, 2, 0, 1, 1, 2)
sync_reset;
check_mem(2034,"100000101","000110010",1,'1'); -- (1, 0, 0, 2, 2, 0, 1, 2, 1)
sync_reset;
check_mem(2035,"100000011","000110100",1,'1'); -- (1, 0, 0, 2, 2, 0, 2, 1, 1)
sync_reset;
check_mem(2036,"100001000","000110000",2,'1'); -- (1, 0, 0, 2, 2, 1, 0, 0, 0)
sync_reset;
check_mem(2037,"100001001","000110000",2,'1'); -- (1, 0, 0, 2, 2, 1, 0, 0, 1)
sync_reset;
check_mem(2038,"100001010","000110000",2,'1'); -- (1, 0, 0, 2, 2, 1, 0, 1, 0)
sync_reset;
check_mem(2039,"100001010","000110001",1,'1'); -- (1, 0, 0, 2, 2, 1, 0, 1, 2)
sync_reset;
check_mem(2040,"100001001","000110010",2,'1'); -- (1, 0, 0, 2, 2, 1, 0, 2, 1)
sync_reset;
check_mem(2041,"100001100","000110000",1,'1'); -- (1, 0, 0, 2, 2, 1, 1, 0, 0)
sync_reset;
check_mem(2042,"100001100","000110001",1,'1'); -- (1, 0, 0, 2, 2, 1, 1, 0, 2)
sync_reset;
check_mem(2043,"100001110","000110001",1,'1'); -- (1, 0, 0, 2, 2, 1, 1, 1, 2)
sync_reset;
check_mem(2044,"100001100","000110010",1,'1'); -- (1, 0, 0, 2, 2, 1, 1, 2, 0)
sync_reset;
check_mem(2045,"100001101","000110010",1,'1'); -- (1, 0, 0, 2, 2, 1, 1, 2, 1)
sync_reset;
check_mem(2046,"100001001","000110100",2,'1'); -- (1, 0, 0, 2, 2, 1, 2, 0, 1)
sync_reset;
check_mem(2047,"100001010","000110100",2,'1'); -- (1, 0, 0, 2, 2, 1, 2, 1, 0)
sync_reset;
check_mem(2048,"100001011","000110100",2,'1'); -- (1, 0, 0, 2, 2, 1, 2, 1, 1)
sync_reset;
check_mem(2049,"101000000","000000001",1,'1'); -- (1, 0, 1, 0, 0, 0, 0, 0, 2)
sync_reset;
check_mem(2050,"101000000","000000010",1,'1'); -- (1, 0, 1, 0, 0, 0, 0, 2, 0)
sync_reset;
check_mem(2051,"101000000","000000011",1,'1'); -- (1, 0, 1, 0, 0, 0, 0, 2, 2)
sync_reset;
check_mem(2052,"101000100","000000011",1,'1'); -- (1, 0, 1, 0, 0, 0, 1, 2, 2)
sync_reset;
check_mem(2053,"101000000","000000100",1,'1'); -- (1, 0, 1, 0, 0, 0, 2, 0, 0)
sync_reset;
check_mem(2054,"101000000","000000101",1,'1'); -- (1, 0, 1, 0, 0, 0, 2, 0, 2)
sync_reset;
check_mem(2055,"101000010","000000101",1,'1'); -- (1, 0, 1, 0, 0, 0, 2, 1, 2)
sync_reset;
check_mem(2056,"101000000","000000110",1,'1'); -- (1, 0, 1, 0, 0, 0, 2, 2, 0)
sync_reset;
check_mem(2057,"101000001","000000110",1,'1'); -- (1, 0, 1, 0, 0, 0, 2, 2, 1)
sync_reset;
check_mem(2058,"101001000","000000011",1,'1'); -- (1, 0, 1, 0, 0, 1, 0, 2, 2)
sync_reset;
check_mem(2059,"101001000","000000101",7,'1'); -- (1, 0, 1, 0, 0, 1, 2, 0, 2)
sync_reset;
check_mem(2060,"101001000","000000110",8,'1'); -- (1, 0, 1, 0, 0, 1, 2, 2, 0)
sync_reset;
check_mem(2061,"101000000","000001000",1,'1'); -- (1, 0, 1, 0, 0, 2, 0, 0, 0)
sync_reset;
check_mem(2062,"101000000","000001001",1,'1'); -- (1, 0, 1, 0, 0, 2, 0, 0, 2)
sync_reset;
check_mem(2063,"101000010","000001001",1,'1'); -- (1, 0, 1, 0, 0, 2, 0, 1, 2)
sync_reset;
check_mem(2064,"101000000","000001010",1,'1'); -- (1, 0, 1, 0, 0, 2, 0, 2, 0)
sync_reset;
check_mem(2065,"101000001","000001010",1,'1'); -- (1, 0, 1, 0, 0, 2, 0, 2, 1)
sync_reset;
check_mem(2066,"101000100","000001001",1,'1'); -- (1, 0, 1, 0, 0, 2, 1, 0, 2)
sync_reset;
check_mem(2067,"101000100","000001010",1,'1'); -- (1, 0, 1, 0, 0, 2, 1, 2, 0)
sync_reset;
check_mem(2068,"101000100","000001011",1,'1'); -- (1, 0, 1, 0, 0, 2, 1, 2, 2)
sync_reset;
check_mem(2069,"101000000","000001100",1,'1'); -- (1, 0, 1, 0, 0, 2, 2, 0, 0)
sync_reset;
check_mem(2070,"101000001","000001100",1,'1'); -- (1, 0, 1, 0, 0, 2, 2, 0, 1)
sync_reset;
check_mem(2071,"101000010","000001100",1,'1'); -- (1, 0, 1, 0, 0, 2, 2, 1, 0)
sync_reset;
check_mem(2072,"101000010","000001101",1,'1'); -- (1, 0, 1, 0, 0, 2, 2, 1, 2)
sync_reset;
check_mem(2073,"101000001","000001110",1,'1'); -- (1, 0, 1, 0, 0, 2, 2, 2, 1)
sync_reset;
check_mem(2074,"101010000","000000011",6,'1'); -- (1, 0, 1, 0, 1, 0, 0, 2, 2)
sync_reset;
check_mem(2075,"101010000","000000101",7,'1'); -- (1, 0, 1, 0, 1, 0, 2, 0, 2)
sync_reset;
check_mem(2076,"101010000","000000110",8,'1'); -- (1, 0, 1, 0, 1, 0, 2, 2, 0)
sync_reset;
check_mem(2077,"101010000","000001001",1,'1'); -- (1, 0, 1, 0, 1, 2, 0, 0, 2)
sync_reset;
check_mem(2078,"101010000","000001010",1,'1'); -- (1, 0, 1, 0, 1, 2, 0, 2, 0)
sync_reset;
check_mem(2079,"101010000","000001011",1,'1'); -- (1, 0, 1, 0, 1, 2, 0, 2, 2)
sync_reset;
check_mem(2080,"101010000","000001100",1,'1'); -- (1, 0, 1, 0, 1, 2, 2, 0, 0)
sync_reset;
check_mem(2081,"101010000","000001101",1,'1'); -- (1, 0, 1, 0, 1, 2, 2, 0, 2)
sync_reset;
check_mem(2082,"101010010","000001101",1,'1'); -- (1, 0, 1, 0, 1, 2, 2, 1, 2)
sync_reset;
check_mem(2083,"101010000","000001110",1,'1'); -- (1, 0, 1, 0, 1, 2, 2, 2, 0)
sync_reset;
check_mem(2084,"101000000","000010000",1,'1'); -- (1, 0, 1, 0, 2, 0, 0, 0, 0)
sync_reset;
check_mem(2085,"101000000","000010001",1,'1'); -- (1, 0, 1, 0, 2, 0, 0, 0, 2)
sync_reset;
check_mem(2086,"101000010","000010001",1,'1'); -- (1, 0, 1, 0, 2, 0, 0, 1, 2)
sync_reset;
check_mem(2087,"101000000","000010010",1,'1'); -- (1, 0, 1, 0, 2, 0, 0, 2, 0)
sync_reset;
check_mem(2088,"101000001","000010010",1,'1'); -- (1, 0, 1, 0, 2, 0, 0, 2, 1)
sync_reset;
check_mem(2089,"101000100","000010001",1,'1'); -- (1, 0, 1, 0, 2, 0, 1, 0, 2)
sync_reset;
check_mem(2090,"101000100","000010010",1,'1'); -- (1, 0, 1, 0, 2, 0, 1, 2, 0)
sync_reset;
check_mem(2091,"101000100","000010011",1,'1'); -- (1, 0, 1, 0, 2, 0, 1, 2, 2)
sync_reset;
check_mem(2092,"101000000","000010100",1,'1'); -- (1, 0, 1, 0, 2, 0, 2, 0, 0)
sync_reset;
check_mem(2093,"101000001","000010100",1,'1'); -- (1, 0, 1, 0, 2, 0, 2, 0, 1)
sync_reset;
check_mem(2094,"101000010","000010100",1,'1'); -- (1, 0, 1, 0, 2, 0, 2, 1, 0)
sync_reset;
check_mem(2095,"101000010","000010101",1,'1'); -- (1, 0, 1, 0, 2, 0, 2, 1, 2)
sync_reset;
check_mem(2096,"101000001","000010110",1,'1'); -- (1, 0, 1, 0, 2, 0, 2, 2, 1)
sync_reset;
check_mem(2097,"101001000","000010001",1,'1'); -- (1, 0, 1, 0, 2, 1, 0, 0, 2)
sync_reset;
check_mem(2098,"101001000","000010010",1,'1'); -- (1, 0, 1, 0, 2, 1, 0, 2, 0)
sync_reset;
check_mem(2099,"101001000","000010011",1,'1'); -- (1, 0, 1, 0, 2, 1, 0, 2, 2)
sync_reset;
check_mem(2100,"101001100","000010011",1,'1'); -- (1, 0, 1, 0, 2, 1, 1, 2, 2)
sync_reset;
check_mem(2101,"101001000","000010100",1,'1'); -- (1, 0, 1, 0, 2, 1, 2, 0, 0)
sync_reset;
check_mem(2102,"101001000","000010101",1,'1'); -- (1, 0, 1, 0, 2, 1, 2, 0, 2)
sync_reset;
check_mem(2103,"101001010","000010101",1,'1'); -- (1, 0, 1, 0, 2, 1, 2, 1, 2)
sync_reset;
check_mem(2104,"101001000","000010110",1,'1'); -- (1, 0, 1, 0, 2, 1, 2, 2, 0)
sync_reset;
check_mem(2105,"101000000","000011000",1,'1'); -- (1, 0, 1, 0, 2, 2, 0, 0, 0)
sync_reset;
check_mem(2106,"101000001","000011000",1,'1'); -- (1, 0, 1, 0, 2, 2, 0, 0, 1)
sync_reset;
check_mem(2107,"101000010","000011000",3,'1'); -- (1, 0, 1, 0, 2, 2, 0, 1, 0)
sync_reset;
check_mem(2108,"101000010","000011001",1,'1'); -- (1, 0, 1, 0, 2, 2, 0, 1, 2)
sync_reset;
check_mem(2109,"101000001","000011010",1,'1'); -- (1, 0, 1, 0, 2, 2, 0, 2, 1)
sync_reset;
check_mem(2110,"101000100","000011000",3,'1'); -- (1, 0, 1, 0, 2, 2, 1, 0, 0)
sync_reset;
check_mem(2111,"101000100","000011001",1,'1'); -- (1, 0, 1, 0, 2, 2, 1, 0, 2)
sync_reset;
check_mem(2112,"101000110","000011001",3,'1'); -- (1, 0, 1, 0, 2, 2, 1, 1, 2)
sync_reset;
check_mem(2113,"101000100","000011010",1,'1'); -- (1, 0, 1, 0, 2, 2, 1, 2, 0)
sync_reset;
check_mem(2114,"101000101","000011010",1,'1'); -- (1, 0, 1, 0, 2, 2, 1, 2, 1)
sync_reset;
check_mem(2115,"101000001","000011100",1,'1'); -- (1, 0, 1, 0, 2, 2, 2, 0, 1)
sync_reset;
check_mem(2116,"101000010","000011100",1,'1'); -- (1, 0, 1, 0, 2, 2, 2, 1, 0)
sync_reset;
check_mem(2117,"101000011","000011100",3,'1'); -- (1, 0, 1, 0, 2, 2, 2, 1, 1)
sync_reset;
check_mem(2118,"101100000","000000011",6,'1'); -- (1, 0, 1, 1, 0, 0, 0, 2, 2)
sync_reset;
check_mem(2119,"101100000","000000101",7,'1'); -- (1, 0, 1, 1, 0, 0, 2, 0, 2)
sync_reset;
check_mem(2120,"101100000","000000110",1,'1'); -- (1, 0, 1, 1, 0, 0, 2, 2, 0)
sync_reset;
check_mem(2121,"101100000","000001001",1,'1'); -- (1, 0, 1, 1, 0, 2, 0, 0, 2)
sync_reset;
check_mem(2122,"101100000","000001010",1,'1'); -- (1, 0, 1, 1, 0, 2, 0, 2, 0)
sync_reset;
check_mem(2123,"101100000","000001011",1,'1'); -- (1, 0, 1, 1, 0, 2, 0, 2, 2)
sync_reset;
check_mem(2124,"101100000","000001100",1,'1'); -- (1, 0, 1, 1, 0, 2, 2, 0, 0)
sync_reset;
check_mem(2125,"101100000","000001101",1,'1'); -- (1, 0, 1, 1, 0, 2, 2, 0, 2)
sync_reset;
check_mem(2126,"101100010","000001101",1,'1'); -- (1, 0, 1, 1, 0, 2, 2, 1, 2)
sync_reset;
check_mem(2127,"101100000","000001110",1,'1'); -- (1, 0, 1, 1, 0, 2, 2, 2, 0)
sync_reset;
check_mem(2128,"101100001","000001110",1,'1'); -- (1, 0, 1, 1, 0, 2, 2, 2, 1)
sync_reset;
check_mem(2129,"101110000","000001011",6,'1'); -- (1, 0, 1, 1, 1, 2, 0, 2, 2)
sync_reset;
check_mem(2130,"101110000","000001101",7,'1'); -- (1, 0, 1, 1, 1, 2, 2, 0, 2)
sync_reset;
check_mem(2131,"101110000","000001110",8,'1'); -- (1, 0, 1, 1, 1, 2, 2, 2, 0)
sync_reset;
check_mem(2132,"101100000","000010001",1,'1'); -- (1, 0, 1, 1, 2, 0, 0, 0, 2)
sync_reset;
check_mem(2133,"101100000","000010010",1,'1'); -- (1, 0, 1, 1, 2, 0, 0, 2, 0)
sync_reset;
check_mem(2134,"101100000","000010011",1,'1'); -- (1, 0, 1, 1, 2, 0, 0, 2, 2)
sync_reset;
check_mem(2135,"101100000","000010100",1,'1'); -- (1, 0, 1, 1, 2, 0, 2, 0, 0)
sync_reset;
check_mem(2136,"101100000","000010101",1,'1'); -- (1, 0, 1, 1, 2, 0, 2, 0, 2)
sync_reset;
check_mem(2137,"101100010","000010101",1,'1'); -- (1, 0, 1, 1, 2, 0, 2, 1, 2)
sync_reset;
check_mem(2138,"101100000","000010110",1,'1'); -- (1, 0, 1, 1, 2, 0, 2, 2, 0)
sync_reset;
check_mem(2139,"101100001","000010110",1,'1'); -- (1, 0, 1, 1, 2, 0, 2, 2, 1)
sync_reset;
check_mem(2140,"101101000","000010011",1,'1'); -- (1, 0, 1, 1, 2, 1, 0, 2, 2)
sync_reset;
check_mem(2141,"101101000","000010101",7,'1'); -- (1, 0, 1, 1, 2, 1, 2, 0, 2)
sync_reset;
check_mem(2142,"101101000","000010110",1,'1'); -- (1, 0, 1, 1, 2, 1, 2, 2, 0)
sync_reset;
check_mem(2143,"101100000","000011000",1,'1'); -- (1, 0, 1, 1, 2, 2, 0, 0, 0)
sync_reset;
check_mem(2144,"101100000","000011001",1,'1'); -- (1, 0, 1, 1, 2, 2, 0, 0, 2)
sync_reset;
check_mem(2145,"101100010","000011001",1,'1'); -- (1, 0, 1, 1, 2, 2, 0, 1, 2)
sync_reset;
check_mem(2146,"101100000","000011010",1,'1'); -- (1, 0, 1, 1, 2, 2, 0, 2, 0)
sync_reset;
check_mem(2147,"101100001","000011010",1,'1'); -- (1, 0, 1, 1, 2, 2, 0, 2, 1)
sync_reset;
check_mem(2148,"101100000","000011100",1,'1'); -- (1, 0, 1, 1, 2, 2, 2, 0, 0)
sync_reset;
check_mem(2149,"101100001","000011100",1,'1'); -- (1, 0, 1, 1, 2, 2, 2, 0, 1)
sync_reset;
check_mem(2150,"101100010","000011100",1,'1'); -- (1, 0, 1, 1, 2, 2, 2, 1, 0)
sync_reset;
check_mem(2151,"101100010","000011101",1,'1'); -- (1, 0, 1, 1, 2, 2, 2, 1, 2)
sync_reset;
check_mem(2152,"101100001","000011110",1,'1'); -- (1, 0, 1, 1, 2, 2, 2, 2, 1)
sync_reset;
check_mem(2153,"101000000","000100000",1,'1'); -- (1, 0, 1, 2, 0, 0, 0, 0, 0)
sync_reset;
check_mem(2154,"101000000","000100001",1,'1'); -- (1, 0, 1, 2, 0, 0, 0, 0, 2)
sync_reset;
check_mem(2155,"101000010","000100001",1,'1'); -- (1, 0, 1, 2, 0, 0, 0, 1, 2)
sync_reset;
check_mem(2156,"101000000","000100010",1,'1'); -- (1, 0, 1, 2, 0, 0, 0, 2, 0)
sync_reset;
check_mem(2157,"101000001","000100010",1,'1'); -- (1, 0, 1, 2, 0, 0, 0, 2, 1)
sync_reset;
check_mem(2158,"101000100","000100001",1,'1'); -- (1, 0, 1, 2, 0, 0, 1, 0, 2)
sync_reset;
check_mem(2159,"101000100","000100010",1,'1'); -- (1, 0, 1, 2, 0, 0, 1, 2, 0)
sync_reset;
check_mem(2160,"101000100","000100011",1,'1'); -- (1, 0, 1, 2, 0, 0, 1, 2, 2)
sync_reset;
check_mem(2161,"101000000","000100100",1,'1'); -- (1, 0, 1, 2, 0, 0, 2, 0, 0)
sync_reset;
check_mem(2162,"101000001","000100100",1,'1'); -- (1, 0, 1, 2, 0, 0, 2, 0, 1)
sync_reset;
check_mem(2163,"101000010","000100100",1,'1'); -- (1, 0, 1, 2, 0, 0, 2, 1, 0)
sync_reset;
check_mem(2164,"101000010","000100101",1,'1'); -- (1, 0, 1, 2, 0, 0, 2, 1, 2)
sync_reset;
check_mem(2165,"101000001","000100110",1,'1'); -- (1, 0, 1, 2, 0, 0, 2, 2, 1)
sync_reset;
check_mem(2166,"101001000","000100001",1,'1'); -- (1, 0, 1, 2, 0, 1, 0, 0, 2)
sync_reset;
check_mem(2167,"101001000","000100010",1,'1'); -- (1, 0, 1, 2, 0, 1, 0, 2, 0)
sync_reset;
check_mem(2168,"101001000","000100011",1,'1'); -- (1, 0, 1, 2, 0, 1, 0, 2, 2)
sync_reset;
check_mem(2169,"101001100","000100011",1,'1'); -- (1, 0, 1, 2, 0, 1, 1, 2, 2)
sync_reset;
check_mem(2170,"101001000","000100100",1,'1'); -- (1, 0, 1, 2, 0, 1, 2, 0, 0)
sync_reset;
check_mem(2171,"101001000","000100101",1,'1'); -- (1, 0, 1, 2, 0, 1, 2, 0, 2)
sync_reset;
check_mem(2172,"101001010","000100101",1,'1'); -- (1, 0, 1, 2, 0, 1, 2, 1, 2)
sync_reset;
check_mem(2173,"101001000","000100110",1,'1'); -- (1, 0, 1, 2, 0, 1, 2, 2, 0)
sync_reset;
check_mem(2174,"101000000","000101000",1,'1'); -- (1, 0, 1, 2, 0, 2, 0, 0, 0)
sync_reset;
check_mem(2175,"101000001","000101000",4,'1'); -- (1, 0, 1, 2, 0, 2, 0, 0, 1)
sync_reset;
check_mem(2176,"101000010","000101000",4,'1'); -- (1, 0, 1, 2, 0, 2, 0, 1, 0)
sync_reset;
check_mem(2177,"101000010","000101001",1,'1'); -- (1, 0, 1, 2, 0, 2, 0, 1, 2)
sync_reset;
check_mem(2178,"101000001","000101010",1,'1'); -- (1, 0, 1, 2, 0, 2, 0, 2, 1)
sync_reset;
check_mem(2179,"101000100","000101000",4,'1'); -- (1, 0, 1, 2, 0, 2, 1, 0, 0)
sync_reset;
check_mem(2180,"101000100","000101001",1,'1'); -- (1, 0, 1, 2, 0, 2, 1, 0, 2)
sync_reset;
check_mem(2181,"101000110","000101001",4,'1'); -- (1, 0, 1, 2, 0, 2, 1, 1, 2)
sync_reset;
check_mem(2182,"101000100","000101010",1,'1'); -- (1, 0, 1, 2, 0, 2, 1, 2, 0)
sync_reset;
check_mem(2183,"101000101","000101010",4,'1'); -- (1, 0, 1, 2, 0, 2, 1, 2, 1)
sync_reset;
check_mem(2184,"101000001","000101100",1,'1'); -- (1, 0, 1, 2, 0, 2, 2, 0, 1)
sync_reset;
check_mem(2185,"101000010","000101100",1,'1'); -- (1, 0, 1, 2, 0, 2, 2, 1, 0)
sync_reset;
check_mem(2186,"101000011","000101100",4,'1'); -- (1, 0, 1, 2, 0, 2, 2, 1, 1)
sync_reset;
check_mem(2187,"101010000","000100001",1,'1'); -- (1, 0, 1, 2, 1, 0, 0, 0, 2)
sync_reset;
check_mem(2188,"101010000","000100010",1,'1'); -- (1, 0, 1, 2, 1, 0, 0, 2, 0)
sync_reset;
check_mem(2189,"101010000","000100011",1,'1'); -- (1, 0, 1, 2, 1, 0, 0, 2, 2)
sync_reset;
check_mem(2190,"101010000","000100100",1,'1'); -- (1, 0, 1, 2, 1, 0, 2, 0, 0)
sync_reset;
check_mem(2191,"101010000","000100101",1,'1'); -- (1, 0, 1, 2, 1, 0, 2, 0, 2)
sync_reset;
check_mem(2192,"101010010","000100101",1,'1'); -- (1, 0, 1, 2, 1, 0, 2, 1, 2)
sync_reset;
check_mem(2193,"101010000","000100110",1,'1'); -- (1, 0, 1, 2, 1, 0, 2, 2, 0)
sync_reset;
check_mem(2194,"101011000","000100011",6,'1'); -- (1, 0, 1, 2, 1, 1, 0, 2, 2)
sync_reset;
check_mem(2195,"101011000","000100101",7,'1'); -- (1, 0, 1, 2, 1, 1, 2, 0, 2)
sync_reset;
check_mem(2196,"101011000","000100110",8,'1'); -- (1, 0, 1, 2, 1, 1, 2, 2, 0)
sync_reset;
check_mem(2197,"101010000","000101000",1,'1'); -- (1, 0, 1, 2, 1, 2, 0, 0, 0)
sync_reset;
check_mem(2198,"101010000","000101001",1,'1'); -- (1, 0, 1, 2, 1, 2, 0, 0, 2)
sync_reset;
check_mem(2199,"101010010","000101001",1,'1'); -- (1, 0, 1, 2, 1, 2, 0, 1, 2)
sync_reset;
check_mem(2200,"101010000","000101010",1,'1'); -- (1, 0, 1, 2, 1, 2, 0, 2, 0)
sync_reset;
check_mem(2201,"101010000","000101100",1,'1'); -- (1, 0, 1, 2, 1, 2, 2, 0, 0)
sync_reset;
check_mem(2202,"101010010","000101100",1,'1'); -- (1, 0, 1, 2, 1, 2, 2, 1, 0)
sync_reset;
check_mem(2203,"101010010","000101101",1,'1'); -- (1, 0, 1, 2, 1, 2, 2, 1, 2)
sync_reset;
check_mem(2204,"101000000","000110000",1,'1'); -- (1, 0, 1, 2, 2, 0, 0, 0, 0)
sync_reset;
check_mem(2205,"101000001","000110000",5,'1'); -- (1, 0, 1, 2, 2, 0, 0, 0, 1)
sync_reset;
check_mem(2206,"101000010","000110000",5,'1'); -- (1, 0, 1, 2, 2, 0, 0, 1, 0)
sync_reset;
check_mem(2207,"101000010","000110001",1,'1'); -- (1, 0, 1, 2, 2, 0, 0, 1, 2)
sync_reset;
check_mem(2208,"101000001","000110010",1,'1'); -- (1, 0, 1, 2, 2, 0, 0, 2, 1)
sync_reset;
check_mem(2209,"101000100","000110000",1,'1'); -- (1, 0, 1, 2, 2, 0, 1, 0, 0)
sync_reset;
check_mem(2210,"101000100","000110001",1,'1'); -- (1, 0, 1, 2, 2, 0, 1, 0, 2)
sync_reset;
check_mem(2211,"101000110","000110001",5,'1'); -- (1, 0, 1, 2, 2, 0, 1, 1, 2)
sync_reset;
check_mem(2212,"101000100","000110010",1,'1'); -- (1, 0, 1, 2, 2, 0, 1, 2, 0)
sync_reset;
check_mem(2213,"101000101","000110010",1,'1'); -- (1, 0, 1, 2, 2, 0, 1, 2, 1)
sync_reset;
check_mem(2214,"101000001","000110100",1,'1'); -- (1, 0, 1, 2, 2, 0, 2, 0, 1)
sync_reset;
check_mem(2215,"101000010","000110100",1,'1'); -- (1, 0, 1, 2, 2, 0, 2, 1, 0)
sync_reset;
check_mem(2216,"101000011","000110100",5,'1'); -- (1, 0, 1, 2, 2, 0, 2, 1, 1)
sync_reset;
check_mem(2217,"101001000","000110000",1,'1'); -- (1, 0, 1, 2, 2, 1, 0, 0, 0)
sync_reset;
check_mem(2218,"101001000","000110001",1,'1'); -- (1, 0, 1, 2, 2, 1, 0, 0, 2)
sync_reset;
check_mem(2219,"101001010","000110001",1,'1'); -- (1, 0, 1, 2, 2, 1, 0, 1, 2)
sync_reset;
check_mem(2220,"101001000","000110010",1,'1'); -- (1, 0, 1, 2, 2, 1, 0, 2, 0)
sync_reset;
check_mem(2221,"101001100","000110001",1,'1'); -- (1, 0, 1, 2, 2, 1, 1, 0, 2)
sync_reset;
check_mem(2222,"101001100","000110010",1,'1'); -- (1, 0, 1, 2, 2, 1, 1, 2, 0)
sync_reset;
check_mem(2223,"101001100","000110011",1,'1'); -- (1, 0, 1, 2, 2, 1, 1, 2, 2)
sync_reset;
check_mem(2224,"101001000","000110100",1,'1'); -- (1, 0, 1, 2, 2, 1, 2, 0, 0)
sync_reset;
check_mem(2225,"101001010","000110100",1,'1'); -- (1, 0, 1, 2, 2, 1, 2, 1, 0)
sync_reset;
check_mem(2226,"101001010","000110101",1,'1'); -- (1, 0, 1, 2, 2, 1, 2, 1, 2)
sync_reset;
check_mem(2227,"100000000","001000000",3,'1'); -- (1, 0, 2, 0, 0, 0, 0, 0, 0)
sync_reset;
check_mem(2228,"100000001","001000000",1,'1'); -- (1, 0, 2, 0, 0, 0, 0, 0, 1)
sync_reset;
check_mem(2229,"100000010","001000000",8,'1'); -- (1, 0, 2, 0, 0, 0, 0, 1, 0)
sync_reset;
check_mem(2230,"100000010","001000001",5,'1'); -- (1, 0, 2, 0, 0, 0, 0, 1, 2)
sync_reset;
check_mem(2231,"100000001","001000010",3,'1'); -- (1, 0, 2, 0, 0, 0, 0, 2, 1)
sync_reset;
check_mem(2232,"100000100","001000000",1,'1'); -- (1, 0, 2, 0, 0, 0, 1, 0, 0)
sync_reset;
check_mem(2233,"100000100","001000001",3,'1'); -- (1, 0, 2, 0, 0, 0, 1, 0, 2)
sync_reset;
check_mem(2234,"100000110","001000001",5,'1'); -- (1, 0, 2, 0, 0, 0, 1, 1, 2)
sync_reset;
check_mem(2235,"100000100","001000010",3,'1'); -- (1, 0, 2, 0, 0, 0, 1, 2, 0)
sync_reset;
check_mem(2236,"100000101","001000010",1,'1'); -- (1, 0, 2, 0, 0, 0, 1, 2, 1)
sync_reset;
check_mem(2237,"100000001","001000100",4,'1'); -- (1, 0, 2, 0, 0, 0, 2, 0, 1)
sync_reset;
check_mem(2238,"100000010","001000100",4,'1'); -- (1, 0, 2, 0, 0, 0, 2, 1, 0)
sync_reset;
check_mem(2239,"100000011","001000100",4,'1'); -- (1, 0, 2, 0, 0, 0, 2, 1, 1)
sync_reset;
check_mem(2240,"100001000","001000000",3,'1'); -- (1, 0, 2, 0, 0, 1, 0, 0, 0)
sync_reset;
check_mem(2241,"100001000","001000001",3,'1'); -- (1, 0, 2, 0, 0, 1, 0, 0, 2)
sync_reset;
check_mem(2242,"100001010","001000001",3,'1'); -- (1, 0, 2, 0, 0, 1, 0, 1, 2)
sync_reset;
check_mem(2243,"100001000","001000010",3,'1'); -- (1, 0, 2, 0, 0, 1, 0, 2, 0)
sync_reset;
check_mem(2244,"100001001","001000010",4,'1'); -- (1, 0, 2, 0, 0, 1, 0, 2, 1)
sync_reset;
check_mem(2245,"100001100","001000001",3,'1'); -- (1, 0, 2, 0, 0, 1, 1, 0, 2)
sync_reset;
check_mem(2246,"100001100","001000010",3,'1'); -- (1, 0, 2, 0, 0, 1, 1, 2, 0)
sync_reset;
check_mem(2247,"100001100","001000011",3,'1'); -- (1, 0, 2, 0, 0, 1, 1, 2, 2)
sync_reset;
check_mem(2248,"100001000","001000100",4,'1'); -- (1, 0, 2, 0, 0, 1, 2, 0, 0)
sync_reset;
check_mem(2249,"100001001","001000100",4,'1'); -- (1, 0, 2, 0, 0, 1, 2, 0, 1)
sync_reset;
check_mem(2250,"100001010","001000100",4,'1'); -- (1, 0, 2, 0, 0, 1, 2, 1, 0)
sync_reset;
check_mem(2251,"100001010","001000101",4,'1'); -- (1, 0, 2, 0, 0, 1, 2, 1, 2)
sync_reset;
check_mem(2252,"100001001","001000110",4,'1'); -- (1, 0, 2, 0, 0, 1, 2, 2, 1)
sync_reset;
check_mem(2253,"100000001","001001000",3,'1'); -- (1, 0, 2, 0, 0, 2, 0, 0, 1)
sync_reset;
check_mem(2254,"100000010","001001000",8,'1'); -- (1, 0, 2, 0, 0, 2, 0, 1, 0)
sync_reset;
check_mem(2255,"100000011","001001000",1,'1'); -- (1, 0, 2, 0, 0, 2, 0, 1, 1)
sync_reset;
check_mem(2256,"100000100","001001000",3,'1'); -- (1, 0, 2, 0, 0, 2, 1, 0, 0)
sync_reset;
check_mem(2257,"100000101","001001000",1,'1'); -- (1, 0, 2, 0, 0, 2, 1, 0, 1)
sync_reset;
check_mem(2258,"100000110","001001000",8,'1'); -- (1, 0, 2, 0, 0, 2, 1, 1, 0)
sync_reset;
check_mem(2259,"100000101","001001010",1,'1'); -- (1, 0, 2, 0, 0, 2, 1, 2, 1)
sync_reset;
check_mem(2260,"100000011","001001100",4,'1'); -- (1, 0, 2, 0, 0, 2, 2, 1, 1)
sync_reset;
check_mem(2261,"100010000","001000000",8,'1'); -- (1, 0, 2, 0, 1, 0, 0, 0, 0)
sync_reset;
check_mem(2262,"100010000","001000001",5,'1'); -- (1, 0, 2, 0, 1, 0, 0, 0, 2)
sync_reset;
check_mem(2263,"100010010","001000001",5,'1'); -- (1, 0, 2, 0, 1, 0, 0, 1, 2)
sync_reset;
check_mem(2264,"100010000","001000010",3,'1'); -- (1, 0, 2, 0, 1, 0, 0, 2, 0)
sync_reset;
check_mem(2265,"100010100","001000001",5,'1'); -- (1, 0, 2, 0, 1, 0, 1, 0, 2)
sync_reset;
check_mem(2266,"100010100","001000010",1,'1'); -- (1, 0, 2, 0, 1, 0, 1, 2, 0)
sync_reset;
check_mem(2267,"100010100","001000011",3,'1'); -- (1, 0, 2, 0, 1, 0, 1, 2, 2)
sync_reset;
check_mem(2268,"100010000","001000100",1,'1'); -- (1, 0, 2, 0, 1, 0, 2, 0, 0)
sync_reset;
check_mem(2269,"100010010","001000100",1,'1'); -- (1, 0, 2, 0, 1, 0, 2, 1, 0)
sync_reset;
check_mem(2270,"100010010","001000101",1,'1'); -- (1, 0, 2, 0, 1, 0, 2, 1, 2)
sync_reset;
check_mem(2271,"100011000","001000001",3,'1'); -- (1, 0, 2, 0, 1, 1, 0, 0, 2)
sync_reset;
check_mem(2272,"100011000","001000010",1,'1'); -- (1, 0, 2, 0, 1, 1, 0, 2, 0)
sync_reset;
check_mem(2273,"100011000","001000011",3,'1'); -- (1, 0, 2, 0, 1, 1, 0, 2, 2)
sync_reset;
check_mem(2274,"100011100","001000011",3,'1'); -- (1, 0, 2, 0, 1, 1, 1, 2, 2)
sync_reset;
check_mem(2275,"100011000","001000100",1,'1'); -- (1, 0, 2, 0, 1, 1, 2, 0, 0)
sync_reset;
check_mem(2276,"100011000","001000101",3,'1'); -- (1, 0, 2, 0, 1, 1, 2, 0, 2)
sync_reset;
check_mem(2277,"100011010","001000101",1,'1'); -- (1, 0, 2, 0, 1, 1, 2, 1, 2)
sync_reset;
check_mem(2278,"100011000","001000110",3,'1'); -- (1, 0, 2, 0, 1, 1, 2, 2, 0)
sync_reset;
check_mem(2279,"100010000","001001000",8,'1'); -- (1, 0, 2, 0, 1, 2, 0, 0, 0)
sync_reset;
check_mem(2280,"100010010","001001000",8,'1'); -- (1, 0, 2, 0, 1, 2, 0, 1, 0)
sync_reset;
check_mem(2281,"100010100","001001000",8,'1'); -- (1, 0, 2, 0, 1, 2, 1, 0, 0)
sync_reset;
check_mem(2282,"100010100","001001010",3,'1'); -- (1, 0, 2, 0, 1, 2, 1, 2, 0)
sync_reset;
check_mem(2283,"100010010","001001100",1,'1'); -- (1, 0, 2, 0, 1, 2, 2, 1, 0)
sync_reset;
check_mem(2284,"100000001","001010000",6,'1'); -- (1, 0, 2, 0, 2, 0, 0, 0, 1)
sync_reset;
check_mem(2285,"100000010","001010000",6,'1'); -- (1, 0, 2, 0, 2, 0, 0, 1, 0)
sync_reset;
check_mem(2286,"100000011","001010000",6,'1'); -- (1, 0, 2, 0, 2, 0, 0, 1, 1)
sync_reset;
check_mem(2287,"100000100","001010000",3,'1'); -- (1, 0, 2, 0, 2, 0, 1, 0, 0)
sync_reset;
check_mem(2288,"100000101","001010000",1,'1'); -- (1, 0, 2, 0, 2, 0, 1, 0, 1)
sync_reset;
check_mem(2289,"100000110","001010000",1,'1'); -- (1, 0, 2, 0, 2, 0, 1, 1, 0)
sync_reset;
check_mem(2290,"100000110","001010001",3,'1'); -- (1, 0, 2, 0, 2, 0, 1, 1, 2)
sync_reset;
check_mem(2291,"100000101","001010010",3,'1'); -- (1, 0, 2, 0, 2, 0, 1, 2, 1)
sync_reset;
check_mem(2292,"100001000","001010000",6,'1'); -- (1, 0, 2, 0, 2, 1, 0, 0, 0)
sync_reset;
check_mem(2293,"100001001","001010000",1,'1'); -- (1, 0, 2, 0, 2, 1, 0, 0, 1)
sync_reset;
check_mem(2294,"100001010","001010000",6,'1'); -- (1, 0, 2, 0, 2, 1, 0, 1, 0)
sync_reset;
check_mem(2295,"100001010","001010001",6,'1'); -- (1, 0, 2, 0, 2, 1, 0, 1, 2)
sync_reset;
check_mem(2296,"100001001","001010010",1,'1'); -- (1, 0, 2, 0, 2, 1, 0, 2, 1)
sync_reset;
check_mem(2297,"100001100","001010000",3,'1'); -- (1, 0, 2, 0, 2, 1, 1, 0, 0)
sync_reset;
check_mem(2298,"100001100","001010001",3,'1'); -- (1, 0, 2, 0, 2, 1, 1, 0, 2)
sync_reset;
check_mem(2299,"100001110","001010001",3,'1'); -- (1, 0, 2, 0, 2, 1, 1, 1, 2)
sync_reset;
check_mem(2300,"100001100","001010010",3,'1'); -- (1, 0, 2, 0, 2, 1, 1, 2, 0)
sync_reset;
check_mem(2301,"100001101","001010010",1,'1'); -- (1, 0, 2, 0, 2, 1, 1, 2, 1)
sync_reset;
check_mem(2302,"100000011","001011000",6,'1'); -- (1, 0, 2, 0, 2, 2, 0, 1, 1)
sync_reset;
check_mem(2303,"100000101","001011000",3,'1'); -- (1, 0, 2, 0, 2, 2, 1, 0, 1)
sync_reset;
check_mem(2304,"100000110","001011000",3,'1'); -- (1, 0, 2, 0, 2, 2, 1, 1, 0)
sync_reset;
check_mem(2305,"100100000","001000000",1,'1'); -- (1, 0, 2, 1, 0, 0, 0, 0, 0)
sync_reset;
check_mem(2306,"100100000","001000001",5,'1'); -- (1, 0, 2, 1, 0, 0, 0, 0, 2)
sync_reset;
check_mem(2307,"100100010","001000001",5,'1'); -- (1, 0, 2, 1, 0, 0, 0, 1, 2)
sync_reset;
check_mem(2308,"100100000","001000010",4,'1'); -- (1, 0, 2, 1, 0, 0, 0, 2, 0)
sync_reset;
check_mem(2309,"100100001","001000010",1,'1'); -- (1, 0, 2, 1, 0, 0, 0, 2, 1)
sync_reset;
check_mem(2310,"100100000","001000100",4,'1'); -- (1, 0, 2, 1, 0, 0, 2, 0, 0)
sync_reset;
check_mem(2311,"100100001","001000100",4,'1'); -- (1, 0, 2, 1, 0, 0, 2, 0, 1)
sync_reset;
check_mem(2312,"100100010","001000100",4,'1'); -- (1, 0, 2, 1, 0, 0, 2, 1, 0)
sync_reset;
check_mem(2313,"100100010","001000101",1,'1'); -- (1, 0, 2, 1, 0, 0, 2, 1, 2)
sync_reset;
check_mem(2314,"100100001","001000110",4,'1'); -- (1, 0, 2, 1, 0, 0, 2, 2, 1)
sync_reset;
check_mem(2315,"100101000","001000001",1,'1'); -- (1, 0, 2, 1, 0, 1, 0, 0, 2)
sync_reset;
check_mem(2316,"100101000","001000010",1,'1'); -- (1, 0, 2, 1, 0, 1, 0, 2, 0)
sync_reset;
check_mem(2317,"100101000","001000011",4,'1'); -- (1, 0, 2, 1, 0, 1, 0, 2, 2)
sync_reset;
check_mem(2318,"100101000","001000100",4,'1'); -- (1, 0, 2, 1, 0, 1, 2, 0, 0)
sync_reset;
check_mem(2319,"100101000","001000101",4,'1'); -- (1, 0, 2, 1, 0, 1, 2, 0, 2)
sync_reset;
check_mem(2320,"100101010","001000101",4,'1'); -- (1, 0, 2, 1, 0, 1, 2, 1, 2)
sync_reset;
check_mem(2321,"100101000","001000110",4,'1'); -- (1, 0, 2, 1, 0, 1, 2, 2, 0)
sync_reset;
check_mem(2322,"100101001","001000110",4,'1'); -- (1, 0, 2, 1, 0, 1, 2, 2, 1)
sync_reset;
check_mem(2323,"100100000","001001000",6,'1'); -- (1, 0, 2, 1, 0, 2, 0, 0, 0)
sync_reset;
check_mem(2324,"100100001","001001000",1,'1'); -- (1, 0, 2, 1, 0, 2, 0, 0, 1)
sync_reset;
check_mem(2325,"100100010","001001000",6,'1'); -- (1, 0, 2, 1, 0, 2, 0, 1, 0)
sync_reset;
check_mem(2326,"100100001","001001010",1,'1'); -- (1, 0, 2, 1, 0, 2, 0, 2, 1)
sync_reset;
check_mem(2327,"100100001","001001100",4,'1'); -- (1, 0, 2, 1, 0, 2, 2, 0, 1)
sync_reset;
check_mem(2328,"100100010","001001100",1,'1'); -- (1, 0, 2, 1, 0, 2, 2, 1, 0)
sync_reset;
check_mem(2329,"100100011","001001100",4,'1'); -- (1, 0, 2, 1, 0, 2, 2, 1, 1)
sync_reset;
check_mem(2330,"100110000","001000001",5,'1'); -- (1, 0, 2, 1, 1, 0, 0, 0, 2)
sync_reset;
check_mem(2331,"100110000","001000010",1,'1'); -- (1, 0, 2, 1, 1, 0, 0, 2, 0)
sync_reset;
check_mem(2332,"100110000","001000011",5,'1'); -- (1, 0, 2, 1, 1, 0, 0, 2, 2)
sync_reset;
check_mem(2333,"100110000","001000100",1,'1'); -- (1, 0, 2, 1, 1, 0, 2, 0, 0)
sync_reset;
check_mem(2334,"100110000","001000101",5,'1'); -- (1, 0, 2, 1, 1, 0, 2, 0, 2)
sync_reset;
check_mem(2335,"100110010","001000101",5,'1'); -- (1, 0, 2, 1, 1, 0, 2, 1, 2)
sync_reset;
check_mem(2336,"100110000","001000110",5,'1'); -- (1, 0, 2, 1, 1, 0, 2, 2, 0)
sync_reset;
check_mem(2337,"100110000","001001000",8,'1'); -- (1, 0, 2, 1, 1, 2, 0, 0, 0)
sync_reset;
check_mem(2338,"100110000","001001010",6,'1'); -- (1, 0, 2, 1, 1, 2, 0, 2, 0)
sync_reset;
check_mem(2339,"100110000","001001100",8,'1'); -- (1, 0, 2, 1, 1, 2, 2, 0, 0)
sync_reset;
check_mem(2340,"100110010","001001100",8,'1'); -- (1, 0, 2, 1, 1, 2, 2, 1, 0)
sync_reset;
check_mem(2341,"100100000","001010000",6,'1'); -- (1, 0, 2, 1, 2, 0, 0, 0, 0)
sync_reset;
check_mem(2342,"100100001","001010000",6,'1'); -- (1, 0, 2, 1, 2, 0, 0, 0, 1)
sync_reset;
check_mem(2343,"100100010","001010000",6,'1'); -- (1, 0, 2, 1, 2, 0, 0, 1, 0)
sync_reset;
check_mem(2344,"100100010","001010001",6,'1'); -- (1, 0, 2, 1, 2, 0, 0, 1, 2)
sync_reset;
check_mem(2345,"100100001","001010010",6,'1'); -- (1, 0, 2, 1, 2, 0, 0, 2, 1)
sync_reset;
check_mem(2346,"100101000","001010000",6,'1'); -- (1, 0, 2, 1, 2, 1, 0, 0, 0)
sync_reset;
check_mem(2347,"100101000","001010001",6,'1'); -- (1, 0, 2, 1, 2, 1, 0, 0, 2)
sync_reset;
check_mem(2348,"100101010","001010001",6,'1'); -- (1, 0, 2, 1, 2, 1, 0, 1, 2)
sync_reset;
check_mem(2349,"100101000","001010010",6,'1'); -- (1, 0, 2, 1, 2, 1, 0, 2, 0)
sync_reset;
check_mem(2350,"100101001","001010010",1,'1'); -- (1, 0, 2, 1, 2, 1, 0, 2, 1)
sync_reset;
check_mem(2351,"100100001","001011000",6,'1'); -- (1, 0, 2, 1, 2, 2, 0, 0, 1)
sync_reset;
check_mem(2352,"100100010","001011000",6,'1'); -- (1, 0, 2, 1, 2, 2, 0, 1, 0)
sync_reset;
check_mem(2353,"100100011","001011000",6,'1'); -- (1, 0, 2, 1, 2, 2, 0, 1, 1)
sync_reset;
check_mem(2354,"100000001","001100000",4,'1'); -- (1, 0, 2, 2, 0, 0, 0, 0, 1)
sync_reset;
check_mem(2355,"100000010","001100000",4,'1'); -- (1, 0, 2, 2, 0, 0, 0, 1, 0)
sync_reset;
check_mem(2356,"100000011","001100000",1,'1'); -- (1, 0, 2, 2, 0, 0, 0, 1, 1)
sync_reset;
check_mem(2357,"100000100","001100000",8,'1'); -- (1, 0, 2, 2, 0, 0, 1, 0, 0)
sync_reset;
check_mem(2358,"100000101","001100000",1,'1'); -- (1, 0, 2, 2, 0, 0, 1, 0, 1)
sync_reset;
check_mem(2359,"100000110","001100000",8,'1'); -- (1, 0, 2, 2, 0, 0, 1, 1, 0)
sync_reset;
check_mem(2360,"100000110","001100001",5,'1'); -- (1, 0, 2, 2, 0, 0, 1, 1, 2)
sync_reset;
check_mem(2361,"100000101","001100010",4,'1'); -- (1, 0, 2, 2, 0, 0, 1, 2, 1)
sync_reset;
check_mem(2362,"100000011","001100100",4,'1'); -- (1, 0, 2, 2, 0, 0, 2, 1, 1)
sync_reset;
check_mem(2363,"100001000","001100000",1,'1'); -- (1, 0, 2, 2, 0, 1, 0, 0, 0)
sync_reset;
check_mem(2364,"100001001","001100000",4,'1'); -- (1, 0, 2, 2, 0, 1, 0, 0, 1)
sync_reset;
check_mem(2365,"100001010","001100000",4,'1'); -- (1, 0, 2, 2, 0, 1, 0, 1, 0)
sync_reset;
check_mem(2366,"100001010","001100001",1,'1'); -- (1, 0, 2, 2, 0, 1, 0, 1, 2)
sync_reset;
check_mem(2367,"100001001","001100010",4,'1'); -- (1, 0, 2, 2, 0, 1, 0, 2, 1)
sync_reset;
check_mem(2368,"100001100","001100000",4,'1'); -- (1, 0, 2, 2, 0, 1, 1, 0, 0)
sync_reset;
check_mem(2369,"100001100","001100001",1,'1'); -- (1, 0, 2, 2, 0, 1, 1, 0, 2)
sync_reset;
check_mem(2370,"100001110","001100001",1,'1'); -- (1, 0, 2, 2, 0, 1, 1, 1, 2)
sync_reset;
check_mem(2371,"100001100","001100010",1,'1'); -- (1, 0, 2, 2, 0, 1, 1, 2, 0)
sync_reset;
check_mem(2372,"100001101","001100010",4,'1'); -- (1, 0, 2, 2, 0, 1, 1, 2, 1)
sync_reset;
check_mem(2373,"100001001","001100100",4,'1'); -- (1, 0, 2, 2, 0, 1, 2, 0, 1)
sync_reset;
check_mem(2374,"100001010","001100100",4,'1'); -- (1, 0, 2, 2, 0, 1, 2, 1, 0)
sync_reset;
check_mem(2375,"100001011","001100100",4,'1'); -- (1, 0, 2, 2, 0, 1, 2, 1, 1)
sync_reset;
check_mem(2376,"100000011","001101000",4,'1'); -- (1, 0, 2, 2, 0, 2, 0, 1, 1)
sync_reset;
check_mem(2377,"100000101","001101000",4,'1'); -- (1, 0, 2, 2, 0, 2, 1, 0, 1)
sync_reset;
check_mem(2378,"100000110","001101000",8,'1'); -- (1, 0, 2, 2, 0, 2, 1, 1, 0)
sync_reset;
check_mem(2379,"100010000","001100000",1,'1'); -- (1, 0, 2, 2, 1, 0, 0, 0, 0)
sync_reset;
check_mem(2380,"100010010","001100000",1,'1'); -- (1, 0, 2, 2, 1, 0, 0, 1, 0)
sync_reset;
check_mem(2381,"100010010","001100001",1,'1'); -- (1, 0, 2, 2, 1, 0, 0, 1, 2)
sync_reset;
check_mem(2382,"100010100","001100000",8,'1'); -- (1, 0, 2, 2, 1, 0, 1, 0, 0)
sync_reset;
check_mem(2383,"100010100","001100001",5,'1'); -- (1, 0, 2, 2, 1, 0, 1, 0, 2)
sync_reset;
check_mem(2384,"100010110","001100001",5,'1'); -- (1, 0, 2, 2, 1, 0, 1, 1, 2)
sync_reset;
check_mem(2385,"100010100","001100010",8,'1'); -- (1, 0, 2, 2, 1, 0, 1, 2, 0)
sync_reset;
check_mem(2386,"100010010","001100100",1,'1'); -- (1, 0, 2, 2, 1, 0, 2, 1, 0)
sync_reset;
check_mem(2387,"100011000","001100000",8,'1'); -- (1, 0, 2, 2, 1, 1, 0, 0, 0)
sync_reset;
check_mem(2388,"100011000","001100001",1,'1'); -- (1, 0, 2, 2, 1, 1, 0, 0, 2)
sync_reset;
check_mem(2389,"100011010","001100001",1,'1'); -- (1, 0, 2, 2, 1, 1, 0, 1, 2)
sync_reset;
check_mem(2390,"100011000","001100010",8,'1'); -- (1, 0, 2, 2, 1, 1, 0, 2, 0)
sync_reset;
check_mem(2391,"100011100","001100001",1,'1'); -- (1, 0, 2, 2, 1, 1, 1, 0, 2)
sync_reset;
check_mem(2392,"100011100","001100010",8,'1'); -- (1, 0, 2, 2, 1, 1, 1, 2, 0)
sync_reset;
check_mem(2393,"100011100","001100011",1,'1'); -- (1, 0, 2, 2, 1, 1, 1, 2, 2)
sync_reset;
check_mem(2394,"100011000","001100100",1,'1'); -- (1, 0, 2, 2, 1, 1, 2, 0, 0)
sync_reset;
check_mem(2395,"100011010","001100100",1,'1'); -- (1, 0, 2, 2, 1, 1, 2, 1, 0)
sync_reset;
check_mem(2396,"100011010","001100101",1,'1'); -- (1, 0, 2, 2, 1, 1, 2, 1, 2)
sync_reset;
check_mem(2397,"100010010","001101000",1,'1'); -- (1, 0, 2, 2, 1, 2, 0, 1, 0)
sync_reset;
check_mem(2398,"100010100","001101000",8,'1'); -- (1, 0, 2, 2, 1, 2, 1, 0, 0)
sync_reset;
check_mem(2399,"100010110","001101000",8,'1'); -- (1, 0, 2, 2, 1, 2, 1, 1, 0)
sync_reset;
check_mem(2400,"100000011","001110000",6,'1'); -- (1, 0, 2, 2, 2, 0, 0, 1, 1)
sync_reset;
check_mem(2401,"100000101","001110000",7,'1'); -- (1, 0, 2, 2, 2, 0, 1, 0, 1)
sync_reset;
check_mem(2402,"100000110","001110000",8,'1'); -- (1, 0, 2, 2, 2, 0, 1, 1, 0)
sync_reset;
check_mem(2403,"100001001","001110000",6,'1'); -- (1, 0, 2, 2, 2, 1, 0, 0, 1)
sync_reset;
check_mem(2404,"100001010","001110000",6,'1'); -- (1, 0, 2, 2, 2, 1, 0, 1, 0)
sync_reset;
check_mem(2405,"100001011","001110000",6,'1'); -- (1, 0, 2, 2, 2, 1, 0, 1, 1)
sync_reset;
check_mem(2406,"100001100","001110000",1,'1'); -- (1, 0, 2, 2, 2, 1, 1, 0, 0)
sync_reset;
check_mem(2407,"100001101","001110000",7,'1'); -- (1, 0, 2, 2, 2, 1, 1, 0, 1)
sync_reset;
check_mem(2408,"100001110","001110000",8,'1'); -- (1, 0, 2, 2, 2, 1, 1, 1, 0)
sync_reset;
check_mem(2409,"100001110","001110001",1,'1'); -- (1, 0, 2, 2, 2, 1, 1, 1, 2)
sync_reset;
check_mem(2410,"100001101","001110010",1,'1'); -- (1, 0, 2, 2, 2, 1, 1, 2, 1)
sync_reset;
check_mem(2411,"110000000","000000001",2,'1'); -- (1, 1, 0, 0, 0, 0, 0, 0, 2)
sync_reset;
check_mem(2412,"110000000","000000010",2,'1'); -- (1, 1, 0, 0, 0, 0, 0, 2, 0)
sync_reset;
check_mem(2413,"110000000","000000011",2,'1'); -- (1, 1, 0, 0, 0, 0, 0, 2, 2)
sync_reset;
check_mem(2414,"110000100","000000011",2,'1'); -- (1, 1, 0, 0, 0, 0, 1, 2, 2)
sync_reset;
check_mem(2415,"110000000","000000100",2,'1'); -- (1, 1, 0, 0, 0, 0, 2, 0, 0)
sync_reset;
check_mem(2416,"110000000","000000101",2,'1'); -- (1, 1, 0, 0, 0, 0, 2, 0, 2)
sync_reset;
check_mem(2417,"110000010","000000101",2,'1'); -- (1, 1, 0, 0, 0, 0, 2, 1, 2)
sync_reset;
check_mem(2418,"110000000","000000110",2,'1'); -- (1, 1, 0, 0, 0, 0, 2, 2, 0)
sync_reset;
check_mem(2419,"110000001","000000110",2,'1'); -- (1, 1, 0, 0, 0, 0, 2, 2, 1)
sync_reset;
check_mem(2420,"110001000","000000011",6,'1'); -- (1, 1, 0, 0, 0, 1, 0, 2, 2)
sync_reset;
check_mem(2421,"110001000","000000101",2,'1'); -- (1, 1, 0, 0, 0, 1, 2, 0, 2)
sync_reset;
check_mem(2422,"110001000","000000110",2,'1'); -- (1, 1, 0, 0, 0, 1, 2, 2, 0)
sync_reset;
check_mem(2423,"110000000","000001000",2,'1'); -- (1, 1, 0, 0, 0, 2, 0, 0, 0)
sync_reset;
check_mem(2424,"110000000","000001001",2,'1'); -- (1, 1, 0, 0, 0, 2, 0, 0, 2)
sync_reset;
check_mem(2425,"110000010","000001001",2,'1'); -- (1, 1, 0, 0, 0, 2, 0, 1, 2)
sync_reset;
check_mem(2426,"110000000","000001010",2,'1'); -- (1, 1, 0, 0, 0, 2, 0, 2, 0)
sync_reset;
check_mem(2427,"110000001","000001010",2,'1'); -- (1, 1, 0, 0, 0, 2, 0, 2, 1)
sync_reset;
check_mem(2428,"110000100","000001001",2,'1'); -- (1, 1, 0, 0, 0, 2, 1, 0, 2)
sync_reset;
check_mem(2429,"110000100","000001010",2,'1'); -- (1, 1, 0, 0, 0, 2, 1, 2, 0)
sync_reset;
check_mem(2430,"110000100","000001011",2,'1'); -- (1, 1, 0, 0, 0, 2, 1, 2, 2)
sync_reset;
check_mem(2431,"110000000","000001100",2,'1'); -- (1, 1, 0, 0, 0, 2, 2, 0, 0)
sync_reset;
check_mem(2432,"110000001","000001100",2,'1'); -- (1, 1, 0, 0, 0, 2, 2, 0, 1)
sync_reset;
check_mem(2433,"110000010","000001100",2,'1'); -- (1, 1, 0, 0, 0, 2, 2, 1, 0)
sync_reset;
check_mem(2434,"110000010","000001101",2,'1'); -- (1, 1, 0, 0, 0, 2, 2, 1, 2)
sync_reset;
check_mem(2435,"110000001","000001110",2,'1'); -- (1, 1, 0, 0, 0, 2, 2, 2, 1)
sync_reset;
check_mem(2436,"110010000","000000011",2,'1'); -- (1, 1, 0, 0, 1, 0, 0, 2, 2)
sync_reset;
check_mem(2437,"110010000","000000101",7,'1'); -- (1, 1, 0, 0, 1, 0, 2, 0, 2)
sync_reset;
check_mem(2438,"110010000","000000110",8,'1'); -- (1, 1, 0, 0, 1, 0, 2, 2, 0)
sync_reset;
check_mem(2439,"110010000","000001001",2,'1'); -- (1, 1, 0, 0, 1, 2, 0, 0, 2)
sync_reset;
check_mem(2440,"110010000","000001010",2,'1'); -- (1, 1, 0, 0, 1, 2, 0, 2, 0)
sync_reset;
check_mem(2441,"110010000","000001011",2,'1'); -- (1, 1, 0, 0, 1, 2, 0, 2, 2)
sync_reset;
check_mem(2442,"110010100","000001011",2,'1'); -- (1, 1, 0, 0, 1, 2, 1, 2, 2)
sync_reset;
check_mem(2443,"110010000","000001100",2,'1'); -- (1, 1, 0, 0, 1, 2, 2, 0, 0)
sync_reset;
check_mem(2444,"110010000","000001101",2,'1'); -- (1, 1, 0, 0, 1, 2, 2, 0, 2)
sync_reset;
check_mem(2445,"110010000","000001110",2,'1'); -- (1, 1, 0, 0, 1, 2, 2, 2, 0)
sync_reset;
check_mem(2446,"110000000","000010000",2,'1'); -- (1, 1, 0, 0, 2, 0, 0, 0, 0)
sync_reset;
check_mem(2447,"110000000","000010001",2,'1'); -- (1, 1, 0, 0, 2, 0, 0, 0, 2)
sync_reset;
check_mem(2448,"110000010","000010001",2,'1'); -- (1, 1, 0, 0, 2, 0, 0, 1, 2)
sync_reset;
check_mem(2449,"110000000","000010010",2,'1'); -- (1, 1, 0, 0, 2, 0, 0, 2, 0)
sync_reset;
check_mem(2450,"110000001","000010010",2,'1'); -- (1, 1, 0, 0, 2, 0, 0, 2, 1)
sync_reset;
check_mem(2451,"110000100","000010001",2,'1'); -- (1, 1, 0, 0, 2, 0, 1, 0, 2)
sync_reset;
check_mem(2452,"110000100","000010010",2,'1'); -- (1, 1, 0, 0, 2, 0, 1, 2, 0)
sync_reset;
check_mem(2453,"110000100","000010011",2,'1'); -- (1, 1, 0, 0, 2, 0, 1, 2, 2)
sync_reset;
check_mem(2454,"110000000","000010100",2,'1'); -- (1, 1, 0, 0, 2, 0, 2, 0, 0)
sync_reset;
check_mem(2455,"110000001","000010100",2,'1'); -- (1, 1, 0, 0, 2, 0, 2, 0, 1)
sync_reset;
check_mem(2456,"110000010","000010100",2,'1'); -- (1, 1, 0, 0, 2, 0, 2, 1, 0)
sync_reset;
check_mem(2457,"110000010","000010101",2,'1'); -- (1, 1, 0, 0, 2, 0, 2, 1, 2)
sync_reset;
check_mem(2458,"110000001","000010110",2,'1'); -- (1, 1, 0, 0, 2, 0, 2, 2, 1)
sync_reset;
check_mem(2459,"110001000","000010001",2,'1'); -- (1, 1, 0, 0, 2, 1, 0, 0, 2)
sync_reset;
check_mem(2460,"110001000","000010010",2,'1'); -- (1, 1, 0, 0, 2, 1, 0, 2, 0)
sync_reset;
check_mem(2461,"110001000","000010011",2,'1'); -- (1, 1, 0, 0, 2, 1, 0, 2, 2)
sync_reset;
check_mem(2462,"110001100","000010011",2,'1'); -- (1, 1, 0, 0, 2, 1, 1, 2, 2)
sync_reset;
check_mem(2463,"110001000","000010100",2,'1'); -- (1, 1, 0, 0, 2, 1, 2, 0, 0)
sync_reset;
check_mem(2464,"110001000","000010101",2,'1'); -- (1, 1, 0, 0, 2, 1, 2, 0, 2)
sync_reset;
check_mem(2465,"110001010","000010101",2,'1'); -- (1, 1, 0, 0, 2, 1, 2, 1, 2)
sync_reset;
check_mem(2466,"110001000","000010110",2,'1'); -- (1, 1, 0, 0, 2, 1, 2, 2, 0)
sync_reset;
check_mem(2467,"110001001","000010110",2,'1'); -- (1, 1, 0, 0, 2, 1, 2, 2, 1)
sync_reset;
check_mem(2468,"110000000","000011000",2,'1'); -- (1, 1, 0, 0, 2, 2, 0, 0, 0)
sync_reset;
check_mem(2469,"110000001","000011000",2,'1'); -- (1, 1, 0, 0, 2, 2, 0, 0, 1)
sync_reset;
check_mem(2470,"110000010","000011000",2,'1'); -- (1, 1, 0, 0, 2, 2, 0, 1, 0)
sync_reset;
check_mem(2471,"110000010","000011001",2,'1'); -- (1, 1, 0, 0, 2, 2, 0, 1, 2)
sync_reset;
check_mem(2472,"110000001","000011010",2,'1'); -- (1, 1, 0, 0, 2, 2, 0, 2, 1)
sync_reset;
check_mem(2473,"110000100","000011000",3,'1'); -- (1, 1, 0, 0, 2, 2, 1, 0, 0)
sync_reset;
check_mem(2474,"110000100","000011001",2,'1'); -- (1, 1, 0, 0, 2, 2, 1, 0, 2)
sync_reset;
check_mem(2475,"110000110","000011001",2,'1'); -- (1, 1, 0, 0, 2, 2, 1, 1, 2)
sync_reset;
check_mem(2476,"110000100","000011010",2,'1'); -- (1, 1, 0, 0, 2, 2, 1, 2, 0)
sync_reset;
check_mem(2477,"110000101","000011010",3,'1'); -- (1, 1, 0, 0, 2, 2, 1, 2, 1)
sync_reset;
check_mem(2478,"110000001","000011100",2,'1'); -- (1, 1, 0, 0, 2, 2, 2, 0, 1)
sync_reset;
check_mem(2479,"110000010","000011100",2,'1'); -- (1, 1, 0, 0, 2, 2, 2, 1, 0)
sync_reset;
check_mem(2480,"110000011","000011100",2,'1'); -- (1, 1, 0, 0, 2, 2, 2, 1, 1)
sync_reset;
check_mem(2481,"110100000","000000011",6,'1'); -- (1, 1, 0, 1, 0, 0, 0, 2, 2)
sync_reset;
check_mem(2482,"110100000","000000101",2,'1'); -- (1, 1, 0, 1, 0, 0, 2, 0, 2)
sync_reset;
check_mem(2483,"110100000","000000110",2,'1'); -- (1, 1, 0, 1, 0, 0, 2, 2, 0)
sync_reset;
check_mem(2484,"110100000","000001001",2,'1'); -- (1, 1, 0, 1, 0, 2, 0, 0, 2)
sync_reset;
check_mem(2485,"110100000","000001010",2,'1'); -- (1, 1, 0, 1, 0, 2, 0, 2, 0)
sync_reset;
check_mem(2486,"110100000","000001011",2,'1'); -- (1, 1, 0, 1, 0, 2, 0, 2, 2)
sync_reset;
check_mem(2487,"110100000","000001100",2,'1'); -- (1, 1, 0, 1, 0, 2, 2, 0, 0)
sync_reset;
check_mem(2488,"110100000","000001101",2,'1'); -- (1, 1, 0, 1, 0, 2, 2, 0, 2)
sync_reset;
check_mem(2489,"110100010","000001101",2,'1'); -- (1, 1, 0, 1, 0, 2, 2, 1, 2)
sync_reset;
check_mem(2490,"110100000","000001110",2,'1'); -- (1, 1, 0, 1, 0, 2, 2, 2, 0)
sync_reset;
check_mem(2491,"110100001","000001110",2,'1'); -- (1, 1, 0, 1, 0, 2, 2, 2, 1)
sync_reset;
check_mem(2492,"110110000","000001011",2,'1'); -- (1, 1, 0, 1, 1, 2, 0, 2, 2)
sync_reset;
check_mem(2493,"110110000","000001101",2,'1'); -- (1, 1, 0, 1, 1, 2, 2, 0, 2)
sync_reset;
check_mem(2494,"110110000","000001110",8,'1'); -- (1, 1, 0, 1, 1, 2, 2, 2, 0)
sync_reset;
check_mem(2495,"110100000","000010001",2,'1'); -- (1, 1, 0, 1, 2, 0, 0, 0, 2)
sync_reset;
check_mem(2496,"110100000","000010010",2,'1'); -- (1, 1, 0, 1, 2, 0, 0, 2, 0)
sync_reset;
check_mem(2497,"110100000","000010011",2,'1'); -- (1, 1, 0, 1, 2, 0, 0, 2, 2)
sync_reset;
check_mem(2498,"110100000","000010100",2,'1'); -- (1, 1, 0, 1, 2, 0, 2, 0, 0)
sync_reset;
check_mem(2499,"110100000","000010101",2,'1'); -- (1, 1, 0, 1, 2, 0, 2, 0, 2)
sync_reset;
check_mem(2500,"110100010","000010101",2,'1'); -- (1, 1, 0, 1, 2, 0, 2, 1, 2)
sync_reset;
check_mem(2501,"110100000","000010110",2,'1'); -- (1, 1, 0, 1, 2, 0, 2, 2, 0)
sync_reset;
check_mem(2502,"110100001","000010110",2,'1'); -- (1, 1, 0, 1, 2, 0, 2, 2, 1)
sync_reset;
check_mem(2503,"110101000","000010011",6,'1'); -- (1, 1, 0, 1, 2, 1, 0, 2, 2)
sync_reset;
check_mem(2504,"110101000","000010101",2,'1'); -- (1, 1, 0, 1, 2, 1, 2, 0, 2)
sync_reset;
check_mem(2505,"110101000","000010110",2,'1'); -- (1, 1, 0, 1, 2, 1, 2, 2, 0)
sync_reset;
check_mem(2506,"110100000","000011000",2,'1'); -- (1, 1, 0, 1, 2, 2, 0, 0, 0)
sync_reset;
check_mem(2507,"110100000","000011001",2,'1'); -- (1, 1, 0, 1, 2, 2, 0, 0, 2)
sync_reset;
check_mem(2508,"110100010","000011001",2,'1'); -- (1, 1, 0, 1, 2, 2, 0, 1, 2)
sync_reset;
check_mem(2509,"110100000","000011010",2,'1'); -- (1, 1, 0, 1, 2, 2, 0, 2, 0)
sync_reset;
check_mem(2510,"110100001","000011010",2,'1'); -- (1, 1, 0, 1, 2, 2, 0, 2, 1)
sync_reset;
check_mem(2511,"110100000","000011100",2,'1'); -- (1, 1, 0, 1, 2, 2, 2, 0, 0)
sync_reset;
check_mem(2512,"110100001","000011100",2,'1'); -- (1, 1, 0, 1, 2, 2, 2, 0, 1)
sync_reset;
check_mem(2513,"110100010","000011100",2,'1'); -- (1, 1, 0, 1, 2, 2, 2, 1, 0)
sync_reset;
check_mem(2514,"110100010","000011101",2,'1'); -- (1, 1, 0, 1, 2, 2, 2, 1, 2)
sync_reset;
check_mem(2515,"110100001","000011110",2,'1'); -- (1, 1, 0, 1, 2, 2, 2, 2, 1)
sync_reset;
check_mem(2516,"110000000","000100000",2,'1'); -- (1, 1, 0, 2, 0, 0, 0, 0, 0)
sync_reset;
check_mem(2517,"110000000","000100001",2,'1'); -- (1, 1, 0, 2, 0, 0, 0, 0, 2)
sync_reset;
check_mem(2518,"110000010","000100001",2,'1'); -- (1, 1, 0, 2, 0, 0, 0, 1, 2)
sync_reset;
check_mem(2519,"110000000","000100010",2,'1'); -- (1, 1, 0, 2, 0, 0, 0, 2, 0)
sync_reset;
check_mem(2520,"110000001","000100010",2,'1'); -- (1, 1, 0, 2, 0, 0, 0, 2, 1)
sync_reset;
check_mem(2521,"110000100","000100001",2,'1'); -- (1, 1, 0, 2, 0, 0, 1, 0, 2)
sync_reset;
check_mem(2522,"110000100","000100010",2,'1'); -- (1, 1, 0, 2, 0, 0, 1, 2, 0)
sync_reset;
check_mem(2523,"110000100","000100011",2,'1'); -- (1, 1, 0, 2, 0, 0, 1, 2, 2)
sync_reset;
check_mem(2524,"110000000","000100100",2,'1'); -- (1, 1, 0, 2, 0, 0, 2, 0, 0)
sync_reset;
check_mem(2525,"110000001","000100100",2,'1'); -- (1, 1, 0, 2, 0, 0, 2, 0, 1)
sync_reset;
check_mem(2526,"110000010","000100100",2,'1'); -- (1, 1, 0, 2, 0, 0, 2, 1, 0)
sync_reset;
check_mem(2527,"110000010","000100101",2,'1'); -- (1, 1, 0, 2, 0, 0, 2, 1, 2)
sync_reset;
check_mem(2528,"110000001","000100110",2,'1'); -- (1, 1, 0, 2, 0, 0, 2, 2, 1)
sync_reset;
check_mem(2529,"110001000","000100001",2,'1'); -- (1, 1, 0, 2, 0, 1, 0, 0, 2)
sync_reset;
check_mem(2530,"110001000","000100010",2,'1'); -- (1, 1, 0, 2, 0, 1, 0, 2, 0)
sync_reset;
check_mem(2531,"110001000","000100011",2,'1'); -- (1, 1, 0, 2, 0, 1, 0, 2, 2)
sync_reset;
check_mem(2532,"110001100","000100011",2,'1'); -- (1, 1, 0, 2, 0, 1, 1, 2, 2)
sync_reset;
check_mem(2533,"110001000","000100100",2,'1'); -- (1, 1, 0, 2, 0, 1, 2, 0, 0)
sync_reset;
check_mem(2534,"110001000","000100101",2,'1'); -- (1, 1, 0, 2, 0, 1, 2, 0, 2)
sync_reset;
check_mem(2535,"110001010","000100101",2,'1'); -- (1, 1, 0, 2, 0, 1, 2, 1, 2)
sync_reset;
check_mem(2536,"110001000","000100110",2,'1'); -- (1, 1, 0, 2, 0, 1, 2, 2, 0)
sync_reset;
check_mem(2537,"110001001","000100110",2,'1'); -- (1, 1, 0, 2, 0, 1, 2, 2, 1)
sync_reset;
check_mem(2538,"110000000","000101000",2,'1'); -- (1, 1, 0, 2, 0, 2, 0, 0, 0)
sync_reset;
check_mem(2539,"110000001","000101000",4,'1'); -- (1, 1, 0, 2, 0, 2, 0, 0, 1)
sync_reset;
check_mem(2540,"110000010","000101000",4,'1'); -- (1, 1, 0, 2, 0, 2, 0, 1, 0)
sync_reset;
check_mem(2541,"110000010","000101001",2,'1'); -- (1, 1, 0, 2, 0, 2, 0, 1, 2)
sync_reset;
check_mem(2542,"110000001","000101010",2,'1'); -- (1, 1, 0, 2, 0, 2, 0, 2, 1)
sync_reset;
check_mem(2543,"110000100","000101000",2,'1'); -- (1, 1, 0, 2, 0, 2, 1, 0, 0)
sync_reset;
check_mem(2544,"110000100","000101001",2,'1'); -- (1, 1, 0, 2, 0, 2, 1, 0, 2)
sync_reset;
check_mem(2545,"110000110","000101001",2,'1'); -- (1, 1, 0, 2, 0, 2, 1, 1, 2)
sync_reset;
check_mem(2546,"110000100","000101010",2,'1'); -- (1, 1, 0, 2, 0, 2, 1, 2, 0)
sync_reset;
check_mem(2547,"110000101","000101010",4,'1'); -- (1, 1, 0, 2, 0, 2, 1, 2, 1)
sync_reset;
check_mem(2548,"110000001","000101100",2,'1'); -- (1, 1, 0, 2, 0, 2, 2, 0, 1)
sync_reset;
check_mem(2549,"110000010","000101100",2,'1'); -- (1, 1, 0, 2, 0, 2, 2, 1, 0)
sync_reset;
check_mem(2550,"110000011","000101100",4,'1'); -- (1, 1, 0, 2, 0, 2, 2, 1, 1)
sync_reset;
check_mem(2551,"110010000","000100001",2,'1'); -- (1, 1, 0, 2, 1, 0, 0, 0, 2)
sync_reset;
check_mem(2552,"110010000","000100010",2,'1'); -- (1, 1, 0, 2, 1, 0, 0, 2, 0)
sync_reset;
check_mem(2553,"110010000","000100011",2,'1'); -- (1, 1, 0, 2, 1, 0, 0, 2, 2)
sync_reset;
check_mem(2554,"110010100","000100011",2,'1'); -- (1, 1, 0, 2, 1, 0, 1, 2, 2)
sync_reset;
check_mem(2555,"110010000","000100100",2,'1'); -- (1, 1, 0, 2, 1, 0, 2, 0, 0)
sync_reset;
check_mem(2556,"110010000","000100101",2,'1'); -- (1, 1, 0, 2, 1, 0, 2, 0, 2)
sync_reset;
check_mem(2557,"110010000","000100110",2,'1'); -- (1, 1, 0, 2, 1, 0, 2, 2, 0)
sync_reset;
check_mem(2558,"110011000","000100011",6,'1'); -- (1, 1, 0, 2, 1, 1, 0, 2, 2)
sync_reset;
check_mem(2559,"110011000","000100101",7,'1'); -- (1, 1, 0, 2, 1, 1, 2, 0, 2)
sync_reset;
check_mem(2560,"110011000","000100110",8,'1'); -- (1, 1, 0, 2, 1, 1, 2, 2, 0)
sync_reset;
check_mem(2561,"110010000","000101000",2,'1'); -- (1, 1, 0, 2, 1, 2, 0, 0, 0)
sync_reset;
check_mem(2562,"110010000","000101001",2,'1'); -- (1, 1, 0, 2, 1, 2, 0, 0, 2)
sync_reset;
check_mem(2563,"110010000","000101010",2,'1'); -- (1, 1, 0, 2, 1, 2, 0, 2, 0)
sync_reset;
check_mem(2564,"110010100","000101001",2,'1'); -- (1, 1, 0, 2, 1, 2, 1, 0, 2)
sync_reset;
check_mem(2565,"110010100","000101010",2,'1'); -- (1, 1, 0, 2, 1, 2, 1, 2, 0)
sync_reset;
check_mem(2566,"110010100","000101011",2,'1'); -- (1, 1, 0, 2, 1, 2, 1, 2, 2)
sync_reset;
check_mem(2567,"110010000","000101100",2,'1'); -- (1, 1, 0, 2, 1, 2, 2, 0, 0)
sync_reset;
check_mem(2568,"110000000","000110000",2,'1'); -- (1, 1, 0, 2, 2, 0, 0, 0, 0)
sync_reset;
check_mem(2569,"110000001","000110000",2,'1'); -- (1, 1, 0, 2, 2, 0, 0, 0, 1)
sync_reset;
check_mem(2570,"110000010","000110000",2,'1'); -- (1, 1, 0, 2, 2, 0, 0, 1, 0)
sync_reset;
check_mem(2571,"110000010","000110001",2,'1'); -- (1, 1, 0, 2, 2, 0, 0, 1, 2)
sync_reset;
check_mem(2572,"110000001","000110010",2,'1'); -- (1, 1, 0, 2, 2, 0, 0, 2, 1)
sync_reset;
check_mem(2573,"110000100","000110000",5,'1'); -- (1, 1, 0, 2, 2, 0, 1, 0, 0)
sync_reset;
check_mem(2574,"110000100","000110001",2,'1'); -- (1, 1, 0, 2, 2, 0, 1, 0, 2)
sync_reset;
check_mem(2575,"110000110","000110001",5,'1'); -- (1, 1, 0, 2, 2, 0, 1, 1, 2)
sync_reset;
check_mem(2576,"110000100","000110010",2,'1'); -- (1, 1, 0, 2, 2, 0, 1, 2, 0)
sync_reset;
check_mem(2577,"110000101","000110010",5,'1'); -- (1, 1, 0, 2, 2, 0, 1, 2, 1)
sync_reset;
check_mem(2578,"110000001","000110100",2,'1'); -- (1, 1, 0, 2, 2, 0, 2, 0, 1)
sync_reset;
check_mem(2579,"110000010","000110100",2,'1'); -- (1, 1, 0, 2, 2, 0, 2, 1, 0)
sync_reset;
check_mem(2580,"110000011","000110100",2,'1'); -- (1, 1, 0, 2, 2, 0, 2, 1, 1)
sync_reset;
check_mem(2581,"110001000","000110000",2,'1'); -- (1, 1, 0, 2, 2, 1, 0, 0, 0)
sync_reset;
check_mem(2582,"110001000","000110001",2,'1'); -- (1, 1, 0, 2, 2, 1, 0, 0, 2)
sync_reset;
check_mem(2583,"110001010","000110001",2,'1'); -- (1, 1, 0, 2, 2, 1, 0, 1, 2)
sync_reset;
check_mem(2584,"110001000","000110010",2,'1'); -- (1, 1, 0, 2, 2, 1, 0, 2, 0)
sync_reset;
check_mem(2585,"110001001","000110010",2,'1'); -- (1, 1, 0, 2, 2, 1, 0, 2, 1)
sync_reset;
check_mem(2586,"110001100","000110001",2,'1'); -- (1, 1, 0, 2, 2, 1, 1, 0, 2)
sync_reset;
check_mem(2587,"110001100","000110010",2,'1'); -- (1, 1, 0, 2, 2, 1, 1, 2, 0)
sync_reset;
check_mem(2588,"110001100","000110011",2,'1'); -- (1, 1, 0, 2, 2, 1, 1, 2, 2)
sync_reset;
check_mem(2589,"110001000","000110100",2,'1'); -- (1, 1, 0, 2, 2, 1, 2, 0, 0)
sync_reset;
check_mem(2590,"110001001","000110100",2,'1'); -- (1, 1, 0, 2, 2, 1, 2, 0, 1)
sync_reset;
check_mem(2591,"110001010","000110100",2,'1'); -- (1, 1, 0, 2, 2, 1, 2, 1, 0)
sync_reset;
check_mem(2592,"110001010","000110101",2,'1'); -- (1, 1, 0, 2, 2, 1, 2, 1, 2)
sync_reset;
check_mem(2593,"110001001","000110110",2,'1'); -- (1, 1, 0, 2, 2, 1, 2, 2, 1)
sync_reset;
check_mem(2594,"110000000","001000000",5,'1'); -- (1, 1, 2, 0, 0, 0, 0, 0, 0)
sync_reset;
check_mem(2595,"110000000","001000001",3,'1'); -- (1, 1, 2, 0, 0, 0, 0, 0, 2)
sync_reset;
check_mem(2596,"110000010","001000001",4,'1'); -- (1, 1, 2, 0, 0, 0, 0, 1, 2)
sync_reset;
check_mem(2597,"110000000","001000010",6,'1'); -- (1, 1, 2, 0, 0, 0, 0, 2, 0)
sync_reset;
check_mem(2598,"110000001","001000010",4,'1'); -- (1, 1, 2, 0, 0, 0, 0, 2, 1)
sync_reset;
check_mem(2599,"110000100","001000001",5,'1'); -- (1, 1, 2, 0, 0, 0, 1, 0, 2)
sync_reset;
check_mem(2600,"110000100","001000010",3,'1'); -- (1, 1, 2, 0, 0, 0, 1, 2, 0)
sync_reset;
check_mem(2601,"110000100","001000011",3,'1'); -- (1, 1, 2, 0, 0, 0, 1, 2, 2)
sync_reset;
check_mem(2602,"110000000","001000100",4,'1'); -- (1, 1, 2, 0, 0, 0, 2, 0, 0)
sync_reset;
check_mem(2603,"110000001","001000100",4,'1'); -- (1, 1, 2, 0, 0, 0, 2, 0, 1)
sync_reset;
check_mem(2604,"110000010","001000100",4,'1'); -- (1, 1, 2, 0, 0, 0, 2, 1, 0)
sync_reset;
check_mem(2605,"110000010","001000101",4,'1'); -- (1, 1, 2, 0, 0, 0, 2, 1, 2)
sync_reset;
check_mem(2606,"110000001","001000110",4,'1'); -- (1, 1, 2, 0, 0, 0, 2, 2, 1)
sync_reset;
check_mem(2607,"110001000","001000001",6,'1'); -- (1, 1, 2, 0, 0, 1, 0, 0, 2)
sync_reset;
check_mem(2608,"110001000","001000010",6,'1'); -- (1, 1, 2, 0, 0, 1, 0, 2, 0)
sync_reset;
check_mem(2609,"110001000","001000011",6,'1'); -- (1, 1, 2, 0, 0, 1, 0, 2, 2)
sync_reset;
check_mem(2610,"110001100","001000011",3,'1'); -- (1, 1, 2, 0, 0, 1, 1, 2, 2)
sync_reset;
check_mem(2611,"110001000","001000100",4,'1'); -- (1, 1, 2, 0, 0, 1, 2, 0, 0)
sync_reset;
check_mem(2612,"110001000","001000101",3,'1'); -- (1, 1, 2, 0, 0, 1, 2, 0, 2)
sync_reset;
check_mem(2613,"110001010","001000101",4,'1'); -- (1, 1, 2, 0, 0, 1, 2, 1, 2)
sync_reset;
check_mem(2614,"110001000","001000110",3,'1'); -- (1, 1, 2, 0, 0, 1, 2, 2, 0)
sync_reset;
check_mem(2615,"110001001","001000110",4,'1'); -- (1, 1, 2, 0, 0, 1, 2, 2, 1)
sync_reset;
check_mem(2616,"110000000","001001000",3,'1'); -- (1, 1, 2, 0, 0, 2, 0, 0, 0)
sync_reset;
check_mem(2617,"110000001","001001000",4,'1'); -- (1, 1, 2, 0, 0, 2, 0, 0, 1)
sync_reset;
check_mem(2618,"110000010","001001000",4,'1'); -- (1, 1, 2, 0, 0, 2, 0, 1, 0)
sync_reset;
check_mem(2619,"110000001","001001010",3,'1'); -- (1, 1, 2, 0, 0, 2, 0, 2, 1)
sync_reset;
check_mem(2620,"110000100","001001000",3,'1'); -- (1, 1, 2, 0, 0, 2, 1, 0, 0)
sync_reset;
check_mem(2621,"110000100","001001010",3,'1'); -- (1, 1, 2, 0, 0, 2, 1, 2, 0)
sync_reset;
check_mem(2622,"110000101","001001010",3,'1'); -- (1, 1, 2, 0, 0, 2, 1, 2, 1)
sync_reset;
check_mem(2623,"110000001","001001100",4,'1'); -- (1, 1, 2, 0, 0, 2, 2, 0, 1)
sync_reset;
check_mem(2624,"110000010","001001100",4,'1'); -- (1, 1, 2, 0, 0, 2, 2, 1, 0)
sync_reset;
check_mem(2625,"110000011","001001100",4,'1'); -- (1, 1, 2, 0, 0, 2, 2, 1, 1)
sync_reset;
check_mem(2626,"110010000","001000001",5,'1'); -- (1, 1, 2, 0, 1, 0, 0, 0, 2)
sync_reset;
check_mem(2627,"110010000","001000010",8,'1'); -- (1, 1, 2, 0, 1, 0, 0, 2, 0)
sync_reset;
check_mem(2628,"110010000","001000011",3,'1'); -- (1, 1, 2, 0, 1, 0, 0, 2, 2)
sync_reset;
check_mem(2629,"110010100","001000011",5,'1'); -- (1, 1, 2, 0, 1, 0, 1, 2, 2)
sync_reset;
check_mem(2630,"110010000","001000100",3,'1'); -- (1, 1, 2, 0, 1, 0, 2, 0, 0)
sync_reset;
check_mem(2631,"110010000","001000101",7,'1'); -- (1, 1, 2, 0, 1, 0, 2, 0, 2)
sync_reset;
check_mem(2632,"110010000","001000110",8,'1'); -- (1, 1, 2, 0, 1, 0, 2, 2, 0)
sync_reset;
check_mem(2633,"110011000","001000011",6,'1'); -- (1, 1, 2, 0, 1, 1, 0, 2, 2)
sync_reset;
check_mem(2634,"110011000","001000101",7,'1'); -- (1, 1, 2, 0, 1, 1, 2, 0, 2)
sync_reset;
check_mem(2635,"110011000","001000110",8,'1'); -- (1, 1, 2, 0, 1, 1, 2, 2, 0)
sync_reset;
check_mem(2636,"110010000","001001000",8,'1'); -- (1, 1, 2, 0, 1, 2, 0, 0, 0)
sync_reset;
check_mem(2637,"110010000","001001010",8,'1'); -- (1, 1, 2, 0, 1, 2, 0, 2, 0)
sync_reset;
check_mem(2638,"110010100","001001010",8,'1'); -- (1, 1, 2, 0, 1, 2, 1, 2, 0)
sync_reset;
check_mem(2639,"110010000","001001100",7,'1'); -- (1, 1, 2, 0, 1, 2, 2, 0, 0)
sync_reset;
check_mem(2640,"110000000","001010000",6,'1'); -- (1, 1, 2, 0, 2, 0, 0, 0, 0)
sync_reset;
check_mem(2641,"110000001","001010000",3,'1'); -- (1, 1, 2, 0, 2, 0, 0, 0, 1)
sync_reset;
check_mem(2642,"110000010","001010000",3,'1'); -- (1, 1, 2, 0, 2, 0, 0, 1, 0)
sync_reset;
check_mem(2643,"110000010","001010001",3,'1'); -- (1, 1, 2, 0, 2, 0, 0, 1, 2)
sync_reset;
check_mem(2644,"110000001","001010010",6,'1'); -- (1, 1, 2, 0, 2, 0, 0, 2, 1)
sync_reset;
check_mem(2645,"110000100","001010000",3,'1'); -- (1, 1, 2, 0, 2, 0, 1, 0, 0)
sync_reset;
check_mem(2646,"110000100","001010001",3,'1'); -- (1, 1, 2, 0, 2, 0, 1, 0, 2)
sync_reset;
check_mem(2647,"110000110","001010001",5,'1'); -- (1, 1, 2, 0, 2, 0, 1, 1, 2)
sync_reset;
check_mem(2648,"110000100","001010010",3,'1'); -- (1, 1, 2, 0, 2, 0, 1, 2, 0)
sync_reset;
check_mem(2649,"110000101","001010010",3,'1'); -- (1, 1, 2, 0, 2, 0, 1, 2, 1)
sync_reset;
check_mem(2650,"110001000","001010000",6,'1'); -- (1, 1, 2, 0, 2, 1, 0, 0, 0)
sync_reset;
check_mem(2651,"110001000","001010001",6,'1'); -- (1, 1, 2, 0, 2, 1, 0, 0, 2)
sync_reset;
check_mem(2652,"110001010","001010001",6,'1'); -- (1, 1, 2, 0, 2, 1, 0, 1, 2)
sync_reset;
check_mem(2653,"110001000","001010010",6,'1'); -- (1, 1, 2, 0, 2, 1, 0, 2, 0)
sync_reset;
check_mem(2654,"110001001","001010010",6,'1'); -- (1, 1, 2, 0, 2, 1, 0, 2, 1)
sync_reset;
check_mem(2655,"110001100","001010001",3,'1'); -- (1, 1, 2, 0, 2, 1, 1, 0, 2)
sync_reset;
check_mem(2656,"110001100","001010010",3,'1'); -- (1, 1, 2, 0, 2, 1, 1, 2, 0)
sync_reset;
check_mem(2657,"110001100","001010011",3,'1'); -- (1, 1, 2, 0, 2, 1, 1, 2, 2)
sync_reset;
check_mem(2658,"110000001","001011000",3,'1'); -- (1, 1, 2, 0, 2, 2, 0, 0, 1)
sync_reset;
check_mem(2659,"110000010","001011000",3,'1'); -- (1, 1, 2, 0, 2, 2, 0, 1, 0)
sync_reset;
check_mem(2660,"110000011","001011000",3,'1'); -- (1, 1, 2, 0, 2, 2, 0, 1, 1)
sync_reset;
check_mem(2661,"110000100","001011000",3,'1'); -- (1, 1, 2, 0, 2, 2, 1, 0, 0)
sync_reset;
check_mem(2662,"110000101","001011000",3,'1'); -- (1, 1, 2, 0, 2, 2, 1, 0, 1)
sync_reset;
check_mem(2663,"110000110","001011000",3,'1'); -- (1, 1, 2, 0, 2, 2, 1, 1, 0)
sync_reset;
check_mem(2664,"110000101","001011010",3,'1'); -- (1, 1, 2, 0, 2, 2, 1, 2, 1)
sync_reset;
check_mem(2665,"110100000","001000001",5,'1'); -- (1, 1, 2, 1, 0, 0, 0, 0, 2)
sync_reset;
check_mem(2666,"110100000","001000010",6,'1'); -- (1, 1, 2, 1, 0, 0, 0, 2, 0)
sync_reset;
check_mem(2667,"110100000","001000011",6,'1'); -- (1, 1, 2, 1, 0, 0, 0, 2, 2)
sync_reset;
check_mem(2668,"110100000","001000100",4,'1'); -- (1, 1, 2, 1, 0, 0, 2, 0, 0)
sync_reset;
check_mem(2669,"110100000","001000101",4,'1'); -- (1, 1, 2, 1, 0, 0, 2, 0, 2)
sync_reset;
check_mem(2670,"110100010","001000101",4,'1'); -- (1, 1, 2, 1, 0, 0, 2, 1, 2)
sync_reset;
check_mem(2671,"110100000","001000110",4,'1'); -- (1, 1, 2, 1, 0, 0, 2, 2, 0)
sync_reset;
check_mem(2672,"110100001","001000110",4,'1'); -- (1, 1, 2, 1, 0, 0, 2, 2, 1)
sync_reset;
check_mem(2673,"110101000","001000011",6,'1'); -- (1, 1, 2, 1, 0, 1, 0, 2, 2)
sync_reset;
check_mem(2674,"110101000","001000101",4,'1'); -- (1, 1, 2, 1, 0, 1, 2, 0, 2)
sync_reset;
check_mem(2675,"110101000","001000110",4,'1'); -- (1, 1, 2, 1, 0, 1, 2, 2, 0)
sync_reset;
check_mem(2676,"110100000","001001000",6,'1'); -- (1, 1, 2, 1, 0, 2, 0, 0, 0)
sync_reset;
check_mem(2677,"110100000","001001010",6,'1'); -- (1, 1, 2, 1, 0, 2, 0, 2, 0)
sync_reset;
check_mem(2678,"110100001","001001010",4,'1'); -- (1, 1, 2, 1, 0, 2, 0, 2, 1)
sync_reset;
check_mem(2679,"110100000","001001100",4,'1'); -- (1, 1, 2, 1, 0, 2, 2, 0, 0)
sync_reset;
check_mem(2680,"110100001","001001100",4,'1'); -- (1, 1, 2, 1, 0, 2, 2, 0, 1)
sync_reset;
check_mem(2681,"110100010","001001100",4,'1'); -- (1, 1, 2, 1, 0, 2, 2, 1, 0)
sync_reset;
check_mem(2682,"110100001","001001110",4,'1'); -- (1, 1, 2, 1, 0, 2, 2, 2, 1)
sync_reset;
check_mem(2683,"110110000","001000011",5,'1'); -- (1, 1, 2, 1, 1, 0, 0, 2, 2)
sync_reset;
check_mem(2684,"110110000","001000101",5,'1'); -- (1, 1, 2, 1, 1, 0, 2, 0, 2)
sync_reset;
check_mem(2685,"110110000","001000110",8,'1'); -- (1, 1, 2, 1, 1, 0, 2, 2, 0)
sync_reset;
check_mem(2686,"110110000","001001010",8,'1'); -- (1, 1, 2, 1, 1, 2, 0, 2, 0)
sync_reset;
check_mem(2687,"110110000","001001100",8,'1'); -- (1, 1, 2, 1, 1, 2, 2, 0, 0)
sync_reset;
check_mem(2688,"110110000","001001110",8,'1'); -- (1, 1, 2, 1, 1, 2, 2, 2, 0)
sync_reset;
check_mem(2689,"110100000","001010000",6,'1'); -- (1, 1, 2, 1, 2, 0, 0, 0, 0)
sync_reset;
check_mem(2690,"110100000","001010001",6,'1'); -- (1, 1, 2, 1, 2, 0, 0, 0, 2)
sync_reset;
check_mem(2691,"110100010","001010001",5,'1'); -- (1, 1, 2, 1, 2, 0, 0, 1, 2)
sync_reset;
check_mem(2692,"110100000","001010010",6,'1'); -- (1, 1, 2, 1, 2, 0, 0, 2, 0)
sync_reset;
check_mem(2693,"110100001","001010010",6,'1'); -- (1, 1, 2, 1, 2, 0, 0, 2, 1)
sync_reset;
check_mem(2694,"110101000","001010001",6,'1'); -- (1, 1, 2, 1, 2, 1, 0, 0, 2)
sync_reset;
check_mem(2695,"110101000","001010010",6,'1'); -- (1, 1, 2, 1, 2, 1, 0, 2, 0)
sync_reset;
check_mem(2696,"110101000","001010011",6,'1'); -- (1, 1, 2, 1, 2, 1, 0, 2, 2)
sync_reset;
check_mem(2697,"110100000","001011000",6,'1'); -- (1, 1, 2, 1, 2, 2, 0, 0, 0)
sync_reset;
check_mem(2698,"110100001","001011000",6,'1'); -- (1, 1, 2, 1, 2, 2, 0, 0, 1)
sync_reset;
check_mem(2699,"110100010","001011000",6,'1'); -- (1, 1, 2, 1, 2, 2, 0, 1, 0)
sync_reset;
check_mem(2700,"110100001","001011010",6,'1'); -- (1, 1, 2, 1, 2, 2, 0, 2, 1)
sync_reset;
check_mem(2701,"110000000","001100000",4,'1'); -- (1, 1, 2, 2, 0, 0, 0, 0, 0)
sync_reset;
check_mem(2702,"110000001","001100000",4,'1'); -- (1, 1, 2, 2, 0, 0, 0, 0, 1)
sync_reset;
check_mem(2703,"110000010","001100000",4,'1'); -- (1, 1, 2, 2, 0, 0, 0, 1, 0)
sync_reset;
check_mem(2704,"110000010","001100001",4,'1'); -- (1, 1, 2, 2, 0, 0, 0, 1, 2)
sync_reset;
check_mem(2705,"110000001","001100010",4,'1'); -- (1, 1, 2, 2, 0, 0, 0, 2, 1)
sync_reset;
check_mem(2706,"110000100","001100000",5,'1'); -- (1, 1, 2, 2, 0, 0, 1, 0, 0)
sync_reset;
check_mem(2707,"110000100","001100001",5,'1'); -- (1, 1, 2, 2, 0, 0, 1, 0, 2)
sync_reset;
check_mem(2708,"110000110","001100001",5,'1'); -- (1, 1, 2, 2, 0, 0, 1, 1, 2)
sync_reset;
check_mem(2709,"110000100","001100010",4,'1'); -- (1, 1, 2, 2, 0, 0, 1, 2, 0)
sync_reset;
check_mem(2710,"110000101","001100010",4,'1'); -- (1, 1, 2, 2, 0, 0, 1, 2, 1)
sync_reset;
check_mem(2711,"110000001","001100100",4,'1'); -- (1, 1, 2, 2, 0, 0, 2, 0, 1)
sync_reset;
check_mem(2712,"110000010","001100100",4,'1'); -- (1, 1, 2, 2, 0, 0, 2, 1, 0)
sync_reset;
check_mem(2713,"110000011","001100100",4,'1'); -- (1, 1, 2, 2, 0, 0, 2, 1, 1)
sync_reset;
check_mem(2714,"110001000","001100000",4,'1'); -- (1, 1, 2, 2, 0, 1, 0, 0, 0)
sync_reset;
check_mem(2715,"110001000","001100001",4,'1'); -- (1, 1, 2, 2, 0, 1, 0, 0, 2)
sync_reset;
check_mem(2716,"110001010","001100001",4,'1'); -- (1, 1, 2, 2, 0, 1, 0, 1, 2)
sync_reset;
check_mem(2717,"110001000","001100010",4,'1'); -- (1, 1, 2, 2, 0, 1, 0, 2, 0)
sync_reset;
check_mem(2718,"110001001","001100010",4,'1'); -- (1, 1, 2, 2, 0, 1, 0, 2, 1)
sync_reset;
check_mem(2719,"110001100","001100001",4,'1'); -- (1, 1, 2, 2, 0, 1, 1, 0, 2)
sync_reset;
check_mem(2720,"110001100","001100010",4,'1'); -- (1, 1, 2, 2, 0, 1, 1, 2, 0)
sync_reset;
check_mem(2721,"110001100","001100011",4,'1'); -- (1, 1, 2, 2, 0, 1, 1, 2, 2)
sync_reset;
check_mem(2722,"110001000","001100100",4,'1'); -- (1, 1, 2, 2, 0, 1, 2, 0, 0)
sync_reset;
check_mem(2723,"110001001","001100100",4,'1'); -- (1, 1, 2, 2, 0, 1, 2, 0, 1)
sync_reset;
check_mem(2724,"110001010","001100100",4,'1'); -- (1, 1, 2, 2, 0, 1, 2, 1, 0)
sync_reset;
check_mem(2725,"110001010","001100101",4,'1'); -- (1, 1, 2, 2, 0, 1, 2, 1, 2)
sync_reset;
check_mem(2726,"110001001","001100110",4,'1'); -- (1, 1, 2, 2, 0, 1, 2, 2, 1)
sync_reset;
check_mem(2727,"110000001","001101000",4,'1'); -- (1, 1, 2, 2, 0, 2, 0, 0, 1)
sync_reset;
check_mem(2728,"110000010","001101000",4,'1'); -- (1, 1, 2, 2, 0, 2, 0, 1, 0)
sync_reset;
check_mem(2729,"110000011","001101000",4,'1'); -- (1, 1, 2, 2, 0, 2, 0, 1, 1)
sync_reset;
check_mem(2730,"110000100","001101000",4,'1'); -- (1, 1, 2, 2, 0, 2, 1, 0, 0)
sync_reset;
check_mem(2731,"110000101","001101000",4,'1'); -- (1, 1, 2, 2, 0, 2, 1, 0, 1)
sync_reset;
check_mem(2732,"110000110","001101000",4,'1'); -- (1, 1, 2, 2, 0, 2, 1, 1, 0)
sync_reset;
check_mem(2733,"110000101","001101010",4,'1'); -- (1, 1, 2, 2, 0, 2, 1, 2, 1)
sync_reset;
check_mem(2734,"110000011","001101100",4,'1'); -- (1, 1, 2, 2, 0, 2, 2, 1, 1)
sync_reset;
check_mem(2735,"110010000","001100000",5,'1'); -- (1, 1, 2, 2, 1, 0, 0, 0, 0)
sync_reset;
check_mem(2736,"110010000","001100001",7,'1'); -- (1, 1, 2, 2, 1, 0, 0, 0, 2)
sync_reset;
check_mem(2737,"110010000","001100010",8,'1'); -- (1, 1, 2, 2, 1, 0, 0, 2, 0)
sync_reset;
check_mem(2738,"110010100","001100001",5,'1'); -- (1, 1, 2, 2, 1, 0, 1, 0, 2)
sync_reset;
check_mem(2739,"110010100","001100010",8,'1'); -- (1, 1, 2, 2, 1, 0, 1, 2, 0)
sync_reset;
check_mem(2740,"110010100","001100011",5,'1'); -- (1, 1, 2, 2, 1, 0, 1, 2, 2)
sync_reset;
check_mem(2741,"110010000","001100100",5,'1'); -- (1, 1, 2, 2, 1, 0, 2, 0, 0)
sync_reset;
check_mem(2742,"110011000","001100001",7,'1'); -- (1, 1, 2, 2, 1, 1, 0, 0, 2)
sync_reset;
check_mem(2743,"110011000","001100010",8,'1'); -- (1, 1, 2, 2, 1, 1, 0, 2, 0)
sync_reset;
check_mem(2744,"110011000","001100011",6,'1'); -- (1, 1, 2, 2, 1, 1, 0, 2, 2)
sync_reset;
check_mem(2745,"110011000","001100100",7,'1'); -- (1, 1, 2, 2, 1, 1, 2, 0, 0)
sync_reset;
check_mem(2746,"110011000","001100101",7,'1'); -- (1, 1, 2, 2, 1, 1, 2, 0, 2)
sync_reset;
check_mem(2747,"110011000","001100110",8,'1'); -- (1, 1, 2, 2, 1, 1, 2, 2, 0)
sync_reset;
check_mem(2748,"110010000","001101000",7,'1'); -- (1, 1, 2, 2, 1, 2, 0, 0, 0)
sync_reset;
check_mem(2749,"110010100","001101000",8,'1'); -- (1, 1, 2, 2, 1, 2, 1, 0, 0)
sync_reset;
check_mem(2750,"110010100","001101010",8,'1'); -- (1, 1, 2, 2, 1, 2, 1, 2, 0)
sync_reset;
check_mem(2751,"110000001","001110000",5,'1'); -- (1, 1, 2, 2, 2, 0, 0, 0, 1)
sync_reset;
check_mem(2752,"110000010","001110000",5,'1'); -- (1, 1, 2, 2, 2, 0, 0, 1, 0)
sync_reset;
check_mem(2753,"110000011","001110000",5,'1'); -- (1, 1, 2, 2, 2, 0, 0, 1, 1)
sync_reset;
check_mem(2754,"110000100","001110000",5,'1'); -- (1, 1, 2, 2, 2, 0, 1, 0, 0)
sync_reset;
check_mem(2755,"110000101","001110000",5,'1'); -- (1, 1, 2, 2, 2, 0, 1, 0, 1)
sync_reset;
check_mem(2756,"110000110","001110000",5,'1'); -- (1, 1, 2, 2, 2, 0, 1, 1, 0)
sync_reset;
check_mem(2757,"110000110","001110001",5,'1'); -- (1, 1, 2, 2, 2, 0, 1, 1, 2)
sync_reset;
check_mem(2758,"110000101","001110010",5,'1'); -- (1, 1, 2, 2, 2, 0, 1, 2, 1)
sync_reset;
check_mem(2759,"110001000","001110000",6,'1'); -- (1, 1, 2, 2, 2, 1, 0, 0, 0)
sync_reset;
check_mem(2760,"110001001","001110000",6,'1'); -- (1, 1, 2, 2, 2, 1, 0, 0, 1)
sync_reset;
check_mem(2761,"110001010","001110000",6,'1'); -- (1, 1, 2, 2, 2, 1, 0, 1, 0)
sync_reset;
check_mem(2762,"110001010","001110001",6,'1'); -- (1, 1, 2, 2, 2, 1, 0, 1, 2)
sync_reset;
check_mem(2763,"110001001","001110010",6,'1'); -- (1, 1, 2, 2, 2, 1, 0, 2, 1)
sync_reset;
check_mem(2764,"110001100","001110000",7,'1'); -- (1, 1, 2, 2, 2, 1, 1, 0, 0)
sync_reset;
check_mem(2765,"110001100","001110001",7,'1'); -- (1, 1, 2, 2, 2, 1, 1, 0, 2)
sync_reset;
check_mem(2766,"110001100","001110010",8,'1'); -- (1, 1, 2, 2, 2, 1, 1, 2, 0)
sync_reset;
check_mem(2767,"100000000","010000000",3,'1'); -- (1, 2, 0, 0, 0, 0, 0, 0, 0)
sync_reset;
check_mem(2768,"100000001","010000000",4,'1'); -- (1, 2, 0, 0, 0, 0, 0, 0, 1)
sync_reset;
check_mem(2769,"100000010","010000000",6,'1'); -- (1, 2, 0, 0, 0, 0, 0, 1, 0)
sync_reset;
check_mem(2770,"100000010","010000001",2,'1'); -- (1, 2, 0, 0, 0, 0, 0, 1, 2)
sync_reset;
check_mem(2771,"100000001","010000010",4,'1'); -- (1, 2, 0, 0, 0, 0, 0, 2, 1)
sync_reset;
check_mem(2772,"100000100","010000000",2,'1'); -- (1, 2, 0, 0, 0, 0, 1, 0, 0)
sync_reset;
check_mem(2773,"100000100","010000001",2,'1'); -- (1, 2, 0, 0, 0, 0, 1, 0, 2)
sync_reset;
check_mem(2774,"100000110","010000001",3,'1'); -- (1, 2, 0, 0, 0, 0, 1, 1, 2)
sync_reset;
check_mem(2775,"100000100","010000010",3,'1'); -- (1, 2, 0, 0, 0, 0, 1, 2, 0)
sync_reset;
check_mem(2776,"100000101","010000010",4,'1'); -- (1, 2, 0, 0, 0, 0, 1, 2, 1)
sync_reset;
check_mem(2777,"100000001","010000100",2,'1'); -- (1, 2, 0, 0, 0, 0, 2, 0, 1)
sync_reset;
check_mem(2778,"100000010","010000100",2,'1'); -- (1, 2, 0, 0, 0, 0, 2, 1, 0)
sync_reset;
check_mem(2779,"100000011","010000100",4,'1'); -- (1, 2, 0, 0, 0, 0, 2, 1, 1)
sync_reset;
check_mem(2780,"100001000","010000000",4,'1'); -- (1, 2, 0, 0, 0, 1, 0, 0, 0)
sync_reset;
check_mem(2781,"100001000","010000001",3,'1'); -- (1, 2, 0, 0, 0, 1, 0, 0, 2)
sync_reset;
check_mem(2782,"100001010","010000001",3,'1'); -- (1, 2, 0, 0, 0, 1, 0, 1, 2)
sync_reset;
check_mem(2783,"100001000","010000010",4,'1'); -- (1, 2, 0, 0, 0, 1, 0, 2, 0)
sync_reset;
check_mem(2784,"100001001","010000010",4,'1'); -- (1, 2, 0, 0, 0, 1, 0, 2, 1)
sync_reset;
check_mem(2785,"100001100","010000001",3,'1'); -- (1, 2, 0, 0, 0, 1, 1, 0, 2)
sync_reset;
check_mem(2786,"100001100","010000010",4,'1'); -- (1, 2, 0, 0, 0, 1, 1, 2, 0)
sync_reset;
check_mem(2787,"100001100","010000011",3,'1'); -- (1, 2, 0, 0, 0, 1, 1, 2, 2)
sync_reset;
check_mem(2788,"100001000","010000100",4,'1'); -- (1, 2, 0, 0, 0, 1, 2, 0, 0)
sync_reset;
check_mem(2789,"100001001","010000100",2,'1'); -- (1, 2, 0, 0, 0, 1, 2, 0, 1)
sync_reset;
check_mem(2790,"100001010","010000100",4,'1'); -- (1, 2, 0, 0, 0, 1, 2, 1, 0)
sync_reset;
check_mem(2791,"100001010","010000101",2,'1'); -- (1, 2, 0, 0, 0, 1, 2, 1, 2)
sync_reset;
check_mem(2792,"100001001","010000110",2,'1'); -- (1, 2, 0, 0, 0, 1, 2, 2, 1)
sync_reset;
check_mem(2793,"100000001","010001000",3,'1'); -- (1, 2, 0, 0, 0, 2, 0, 0, 1)
sync_reset;
check_mem(2794,"100000010","010001000",6,'1'); -- (1, 2, 0, 0, 0, 2, 0, 1, 0)
sync_reset;
check_mem(2795,"100000011","010001000",2,'1'); -- (1, 2, 0, 0, 0, 2, 0, 1, 1)
sync_reset;
check_mem(2796,"100000100","010001000",2,'1'); -- (1, 2, 0, 0, 0, 2, 1, 0, 0)
sync_reset;
check_mem(2797,"100000101","010001000",2,'1'); -- (1, 2, 0, 0, 0, 2, 1, 0, 1)
sync_reset;
check_mem(2798,"100000110","010001000",2,'1'); -- (1, 2, 0, 0, 0, 2, 1, 1, 0)
sync_reset;
check_mem(2799,"100000110","010001001",2,'1'); -- (1, 2, 0, 0, 0, 2, 1, 1, 2)
sync_reset;
check_mem(2800,"100000101","010001010",3,'1'); -- (1, 2, 0, 0, 0, 2, 1, 2, 1)
sync_reset;
check_mem(2801,"100000011","010001100",4,'1'); -- (1, 2, 0, 0, 0, 2, 2, 1, 1)
sync_reset;
check_mem(2802,"100010000","010000000",2,'1'); -- (1, 2, 0, 0, 1, 0, 0, 0, 0)
sync_reset;
check_mem(2803,"100010000","010000001",3,'1'); -- (1, 2, 0, 0, 1, 0, 0, 0, 2)
sync_reset;
check_mem(2804,"100010010","010000001",2,'1'); -- (1, 2, 0, 0, 1, 0, 0, 1, 2)
sync_reset;
check_mem(2805,"100010000","010000010",2,'1'); -- (1, 2, 0, 0, 1, 0, 0, 2, 0)
sync_reset;
check_mem(2806,"100010100","010000001",2,'1'); -- (1, 2, 0, 0, 1, 0, 1, 0, 2)
sync_reset;
check_mem(2807,"100010100","010000010",2,'1'); -- (1, 2, 0, 0, 1, 0, 1, 2, 0)
sync_reset;
check_mem(2808,"100010100","010000011",2,'1'); -- (1, 2, 0, 0, 1, 0, 1, 2, 2)
sync_reset;
check_mem(2809,"100010000","010000100",3,'1'); -- (1, 2, 0, 0, 1, 0, 2, 0, 0)
sync_reset;
check_mem(2810,"100010010","010000100",8,'1'); -- (1, 2, 0, 0, 1, 0, 2, 1, 0)
sync_reset;
check_mem(2811,"100010010","010000101",2,'1'); -- (1, 2, 0, 0, 1, 0, 2, 1, 2)
sync_reset;
check_mem(2812,"100011000","010000001",3,'1'); -- (1, 2, 0, 0, 1, 1, 0, 0, 2)
sync_reset;
check_mem(2813,"100011000","010000010",2,'1'); -- (1, 2, 0, 0, 1, 1, 0, 2, 0)
sync_reset;
check_mem(2814,"100011000","010000011",3,'1'); -- (1, 2, 0, 0, 1, 1, 0, 2, 2)
sync_reset;
check_mem(2815,"100011100","010000011",2,'1'); -- (1, 2, 0, 0, 1, 1, 1, 2, 2)
sync_reset;
check_mem(2816,"100011000","010000100",2,'1'); -- (1, 2, 0, 0, 1, 1, 2, 0, 0)
sync_reset;
check_mem(2817,"100011000","010000101",3,'1'); -- (1, 2, 0, 0, 1, 1, 2, 0, 2)
sync_reset;
check_mem(2818,"100011010","010000101",3,'1'); -- (1, 2, 0, 0, 1, 1, 2, 1, 2)
sync_reset;
check_mem(2819,"100011000","010000110",3,'1'); -- (1, 2, 0, 0, 1, 1, 2, 2, 0)
sync_reset;
check_mem(2820,"100010000","010001000",2,'1'); -- (1, 2, 0, 0, 1, 2, 0, 0, 0)
sync_reset;
check_mem(2821,"100010010","010001000",8,'1'); -- (1, 2, 0, 0, 1, 2, 0, 1, 0)
sync_reset;
check_mem(2822,"100010010","010001001",2,'1'); -- (1, 2, 0, 0, 1, 2, 0, 1, 2)
sync_reset;
check_mem(2823,"100010100","010001000",2,'1'); -- (1, 2, 0, 0, 1, 2, 1, 0, 0)
sync_reset;
check_mem(2824,"100010100","010001001",2,'1'); -- (1, 2, 0, 0, 1, 2, 1, 0, 2)
sync_reset;
check_mem(2825,"100010110","010001001",2,'1'); -- (1, 2, 0, 0, 1, 2, 1, 1, 2)
sync_reset;
check_mem(2826,"100010100","010001010",2,'1'); -- (1, 2, 0, 0, 1, 2, 1, 2, 0)
sync_reset;
check_mem(2827,"100010010","010001100",8,'1'); -- (1, 2, 0, 0, 1, 2, 2, 1, 0)
sync_reset;
check_mem(2828,"100000001","010010000",7,'1'); -- (1, 2, 0, 0, 2, 0, 0, 0, 1)
sync_reset;
check_mem(2829,"100000010","010010000",6,'1'); -- (1, 2, 0, 0, 2, 0, 0, 1, 0)
sync_reset;
check_mem(2830,"100000011","010010000",6,'1'); -- (1, 2, 0, 0, 2, 0, 0, 1, 1)
sync_reset;
check_mem(2831,"100000100","010010000",3,'1'); -- (1, 2, 0, 0, 2, 0, 1, 0, 0)
sync_reset;
check_mem(2832,"100000101","010010000",7,'1'); -- (1, 2, 0, 0, 2, 0, 1, 0, 1)
sync_reset;
check_mem(2833,"100000110","010010000",2,'1'); -- (1, 2, 0, 0, 2, 0, 1, 1, 0)
sync_reset;
check_mem(2834,"100000110","010010001",3,'1'); -- (1, 2, 0, 0, 2, 0, 1, 1, 2)
sync_reset;
check_mem(2835,"100000011","010010100",2,'1'); -- (1, 2, 0, 0, 2, 0, 2, 1, 1)
sync_reset;
check_mem(2836,"100001000","010010000",7,'1'); -- (1, 2, 0, 0, 2, 1, 0, 0, 0)
sync_reset;
check_mem(2837,"100001001","010010000",2,'1'); -- (1, 2, 0, 0, 2, 1, 0, 0, 1)
sync_reset;
check_mem(2838,"100001010","010010000",6,'1'); -- (1, 2, 0, 0, 2, 1, 0, 1, 0)
sync_reset;
check_mem(2839,"100001010","010010001",2,'1'); -- (1, 2, 0, 0, 2, 1, 0, 1, 2)
sync_reset;
check_mem(2840,"100001100","010010000",7,'1'); -- (1, 2, 0, 0, 2, 1, 1, 0, 0)
sync_reset;
check_mem(2841,"100001100","010010001",3,'1'); -- (1, 2, 0, 0, 2, 1, 1, 0, 2)
sync_reset;
check_mem(2842,"100001110","010010001",3,'1'); -- (1, 2, 0, 0, 2, 1, 1, 1, 2)
sync_reset;
check_mem(2843,"100001001","010010100",2,'1'); -- (1, 2, 0, 0, 2, 1, 2, 0, 1)
sync_reset;
check_mem(2844,"100001010","010010100",2,'1'); -- (1, 2, 0, 0, 2, 1, 2, 1, 0)
sync_reset;
check_mem(2845,"100001011","010010100",2,'1'); -- (1, 2, 0, 0, 2, 1, 2, 1, 1)
sync_reset;
check_mem(2846,"100000011","010011000",6,'1'); -- (1, 2, 0, 0, 2, 2, 0, 1, 1)
sync_reset;
check_mem(2847,"100000101","010011000",3,'1'); -- (1, 2, 0, 0, 2, 2, 1, 0, 1)
sync_reset;
check_mem(2848,"100000110","010011000",3,'1'); -- (1, 2, 0, 0, 2, 2, 1, 1, 0)
sync_reset;
check_mem(2849,"100100000","010000000",2,'1'); -- (1, 2, 0, 1, 0, 0, 0, 0, 0)
sync_reset;
check_mem(2850,"100100000","010000001",4,'1'); -- (1, 2, 0, 1, 0, 0, 0, 0, 2)
sync_reset;
check_mem(2851,"100100010","010000001",6,'1'); -- (1, 2, 0, 1, 0, 0, 0, 1, 2)
sync_reset;
check_mem(2852,"100100000","010000010",4,'1'); -- (1, 2, 0, 1, 0, 0, 0, 2, 0)
sync_reset;
check_mem(2853,"100100001","010000010",4,'1'); -- (1, 2, 0, 1, 0, 0, 0, 2, 1)
sync_reset;
check_mem(2854,"100100000","010000100",4,'1'); -- (1, 2, 0, 1, 0, 0, 2, 0, 0)
sync_reset;
check_mem(2855,"100100001","010000100",4,'1'); -- (1, 2, 0, 1, 0, 0, 2, 0, 1)
sync_reset;
check_mem(2856,"100100010","010000100",4,'1'); -- (1, 2, 0, 1, 0, 0, 2, 1, 0)
sync_reset;
check_mem(2857,"100100010","010000101",2,'1'); -- (1, 2, 0, 1, 0, 0, 2, 1, 2)
sync_reset;
check_mem(2858,"100100001","010000110",4,'1'); -- (1, 2, 0, 1, 0, 0, 2, 2, 1)
sync_reset;
check_mem(2859,"100101000","010000001",2,'1'); -- (1, 2, 0, 1, 0, 1, 0, 0, 2)
sync_reset;
check_mem(2860,"100101000","010000010",4,'1'); -- (1, 2, 0, 1, 0, 1, 0, 2, 0)
sync_reset;
check_mem(2861,"100101000","010000011",4,'1'); -- (1, 2, 0, 1, 0, 1, 0, 2, 2)
sync_reset;
check_mem(2862,"100101000","010000100",4,'1'); -- (1, 2, 0, 1, 0, 1, 2, 0, 0)
sync_reset;
check_mem(2863,"100101000","010000101",4,'1'); -- (1, 2, 0, 1, 0, 1, 2, 0, 2)
sync_reset;
check_mem(2864,"100101010","010000101",4,'1'); -- (1, 2, 0, 1, 0, 1, 2, 1, 2)
sync_reset;
check_mem(2865,"100101000","010000110",4,'1'); -- (1, 2, 0, 1, 0, 1, 2, 2, 0)
sync_reset;
check_mem(2866,"100101001","010000110",4,'1'); -- (1, 2, 0, 1, 0, 1, 2, 2, 1)
sync_reset;
check_mem(2867,"100100000","010001000",4,'1'); -- (1, 2, 0, 1, 0, 2, 0, 0, 0)
sync_reset;
check_mem(2868,"100100001","010001000",2,'1'); -- (1, 2, 0, 1, 0, 2, 0, 0, 1)
sync_reset;
check_mem(2869,"100100010","010001000",6,'1'); -- (1, 2, 0, 1, 0, 2, 0, 1, 0)
sync_reset;
check_mem(2870,"100100010","010001001",6,'1'); -- (1, 2, 0, 1, 0, 2, 0, 1, 2)
sync_reset;
check_mem(2871,"100100001","010001010",4,'1'); -- (1, 2, 0, 1, 0, 2, 0, 2, 1)
sync_reset;
check_mem(2872,"100100001","010001100",4,'1'); -- (1, 2, 0, 1, 0, 2, 2, 0, 1)
sync_reset;
check_mem(2873,"100100010","010001100",2,'1'); -- (1, 2, 0, 1, 0, 2, 2, 1, 0)
sync_reset;
check_mem(2874,"100100011","010001100",4,'1'); -- (1, 2, 0, 1, 0, 2, 2, 1, 1)
sync_reset;
check_mem(2875,"100110000","010000001",2,'1'); -- (1, 2, 0, 1, 1, 0, 0, 0, 2)
sync_reset;
check_mem(2876,"100110000","010000010",2,'1'); -- (1, 2, 0, 1, 1, 0, 0, 2, 0)
sync_reset;
check_mem(2877,"100110000","010000011",5,'1'); -- (1, 2, 0, 1, 1, 0, 0, 2, 2)
sync_reset;
check_mem(2878,"100110000","010000100",2,'1'); -- (1, 2, 0, 1, 1, 0, 2, 0, 0)
sync_reset;
check_mem(2879,"100110000","010000101",5,'1'); -- (1, 2, 0, 1, 1, 0, 2, 0, 2)
sync_reset;
check_mem(2880,"100110010","010000101",5,'1'); -- (1, 2, 0, 1, 1, 0, 2, 1, 2)
sync_reset;
check_mem(2881,"100110000","010000110",5,'1'); -- (1, 2, 0, 1, 1, 0, 2, 2, 0)
sync_reset;
check_mem(2882,"100110000","010001000",2,'1'); -- (1, 2, 0, 1, 1, 2, 0, 0, 0)
sync_reset;
check_mem(2883,"100110000","010001001",6,'1'); -- (1, 2, 0, 1, 1, 2, 0, 0, 2)
sync_reset;
check_mem(2884,"100110010","010001001",2,'1'); -- (1, 2, 0, 1, 1, 2, 0, 1, 2)
sync_reset;
check_mem(2885,"100110000","010001010",2,'1'); -- (1, 2, 0, 1, 1, 2, 0, 2, 0)
sync_reset;
check_mem(2886,"100110000","010001100",8,'1'); -- (1, 2, 0, 1, 1, 2, 2, 0, 0)
sync_reset;
check_mem(2887,"100110010","010001100",8,'1'); -- (1, 2, 0, 1, 1, 2, 2, 1, 0)
sync_reset;
check_mem(2888,"100110010","010001101",2,'1'); -- (1, 2, 0, 1, 1, 2, 2, 1, 2)
sync_reset;
check_mem(2889,"100100000","010010000",6,'1'); -- (1, 2, 0, 1, 2, 0, 0, 0, 0)
sync_reset;
check_mem(2890,"100100001","010010000",6,'1'); -- (1, 2, 0, 1, 2, 0, 0, 0, 1)
sync_reset;
check_mem(2891,"100100010","010010000",6,'1'); -- (1, 2, 0, 1, 2, 0, 0, 1, 0)
sync_reset;
check_mem(2892,"100100010","010010001",6,'1'); -- (1, 2, 0, 1, 2, 0, 0, 1, 2)
sync_reset;
check_mem(2893,"100100001","010010100",2,'1'); -- (1, 2, 0, 1, 2, 0, 2, 0, 1)
sync_reset;
check_mem(2894,"100100010","010010100",2,'1'); -- (1, 2, 0, 1, 2, 0, 2, 1, 0)
sync_reset;
check_mem(2895,"100100011","010010100",2,'1'); -- (1, 2, 0, 1, 2, 0, 2, 1, 1)
sync_reset;
check_mem(2896,"100101000","010010000",6,'1'); -- (1, 2, 0, 1, 2, 1, 0, 0, 0)
sync_reset;
check_mem(2897,"100101000","010010001",6,'1'); -- (1, 2, 0, 1, 2, 1, 0, 0, 2)
sync_reset;
check_mem(2898,"100101010","010010001",6,'1'); -- (1, 2, 0, 1, 2, 1, 0, 1, 2)
sync_reset;
check_mem(2899,"100101000","010010100",2,'1'); -- (1, 2, 0, 1, 2, 1, 2, 0, 0)
sync_reset;
check_mem(2900,"100101001","010010100",2,'1'); -- (1, 2, 0, 1, 2, 1, 2, 0, 1)
sync_reset;
check_mem(2901,"100101010","010010100",2,'1'); -- (1, 2, 0, 1, 2, 1, 2, 1, 0)
sync_reset;
check_mem(2902,"100101010","010010101",2,'1'); -- (1, 2, 0, 1, 2, 1, 2, 1, 2)
sync_reset;
check_mem(2903,"100100001","010011000",6,'1'); -- (1, 2, 0, 1, 2, 2, 0, 0, 1)
sync_reset;
check_mem(2904,"100100010","010011000",6,'1'); -- (1, 2, 0, 1, 2, 2, 0, 1, 0)
sync_reset;
check_mem(2905,"100100011","010011000",6,'1'); -- (1, 2, 0, 1, 2, 2, 0, 1, 1)
sync_reset;
check_mem(2906,"100100011","010011100",2,'1'); -- (1, 2, 0, 1, 2, 2, 2, 1, 1)
sync_reset;
check_mem(2907,"100000001","010100000",2,'1'); -- (1, 2, 0, 2, 0, 0, 0, 0, 1)
sync_reset;
check_mem(2908,"100000010","010100000",8,'1'); -- (1, 2, 0, 2, 0, 0, 0, 1, 0)
sync_reset;
check_mem(2909,"100000011","010100000",2,'1'); -- (1, 2, 0, 2, 0, 0, 0, 1, 1)
sync_reset;
check_mem(2910,"100000100","010100000",4,'1'); -- (1, 2, 0, 2, 0, 0, 1, 0, 0)
sync_reset;
check_mem(2911,"100000101","010100000",2,'1'); -- (1, 2, 0, 2, 0, 0, 1, 0, 1)
sync_reset;
check_mem(2912,"100000110","010100000",8,'1'); -- (1, 2, 0, 2, 0, 0, 1, 1, 0)
sync_reset;
check_mem(2913,"100000110","010100001",2,'1'); -- (1, 2, 0, 2, 0, 0, 1, 1, 2)
sync_reset;
check_mem(2914,"100000101","010100010",4,'1'); -- (1, 2, 0, 2, 0, 0, 1, 2, 1)
sync_reset;
check_mem(2915,"100000011","010100100",2,'1'); -- (1, 2, 0, 2, 0, 0, 2, 1, 1)
sync_reset;
check_mem(2916,"100001000","010100000",8,'1'); -- (1, 2, 0, 2, 0, 1, 0, 0, 0)
sync_reset;
check_mem(2917,"100001001","010100000",2,'1'); -- (1, 2, 0, 2, 0, 1, 0, 0, 1)
sync_reset;
check_mem(2918,"100001010","010100000",8,'1'); -- (1, 2, 0, 2, 0, 1, 0, 1, 0)
sync_reset;
check_mem(2919,"100001010","010100001",2,'1'); -- (1, 2, 0, 2, 0, 1, 0, 1, 2)
sync_reset;
check_mem(2920,"100001001","010100010",2,'1'); -- (1, 2, 0, 2, 0, 1, 0, 2, 1)
sync_reset;
check_mem(2921,"100001100","010100000",4,'1'); -- (1, 2, 0, 2, 0, 1, 1, 0, 0)
sync_reset;
check_mem(2922,"100001100","010100001",2,'1'); -- (1, 2, 0, 2, 0, 1, 1, 0, 2)
sync_reset;
check_mem(2923,"100001110","010100001",2,'1'); -- (1, 2, 0, 2, 0, 1, 1, 1, 2)
sync_reset;
check_mem(2924,"100001100","010100010",4,'1'); -- (1, 2, 0, 2, 0, 1, 1, 2, 0)
sync_reset;
check_mem(2925,"100001101","010100010",4,'1'); -- (1, 2, 0, 2, 0, 1, 1, 2, 1)
sync_reset;
check_mem(2926,"100001001","010100100",2,'1'); -- (1, 2, 0, 2, 0, 1, 2, 0, 1)
sync_reset;
check_mem(2927,"100001010","010100100",8,'1'); -- (1, 2, 0, 2, 0, 1, 2, 1, 0)
sync_reset;
check_mem(2928,"100001011","010100100",2,'1'); -- (1, 2, 0, 2, 0, 1, 2, 1, 1)
sync_reset;
check_mem(2929,"100000011","010101000",4,'1'); -- (1, 2, 0, 2, 0, 2, 0, 1, 1)
sync_reset;
check_mem(2930,"100000101","010101000",4,'1'); -- (1, 2, 0, 2, 0, 2, 1, 0, 1)
sync_reset;
check_mem(2931,"100000110","010101000",4,'1'); -- (1, 2, 0, 2, 0, 2, 1, 1, 0)
sync_reset;
check_mem(2932,"100010000","010100000",2,'1'); -- (1, 2, 0, 2, 1, 0, 0, 0, 0)
sync_reset;
check_mem(2933,"100010010","010100000",8,'1'); -- (1, 2, 0, 2, 1, 0, 0, 1, 0)
sync_reset;
check_mem(2934,"100010010","010100001",2,'1'); -- (1, 2, 0, 2, 1, 0, 0, 1, 2)
sync_reset;
check_mem(2935,"100010100","010100000",2,'1'); -- (1, 2, 0, 2, 1, 0, 1, 0, 0)
sync_reset;
check_mem(2936,"100010100","010100001",2,'1'); -- (1, 2, 0, 2, 1, 0, 1, 0, 2)
sync_reset;
check_mem(2937,"100010110","010100001",2,'1'); -- (1, 2, 0, 2, 1, 0, 1, 1, 2)
sync_reset;
check_mem(2938,"100010100","010100010",2,'1'); -- (1, 2, 0, 2, 1, 0, 1, 2, 0)
sync_reset;
check_mem(2939,"100010010","010100100",8,'1'); -- (1, 2, 0, 2, 1, 0, 2, 1, 0)
sync_reset;
check_mem(2940,"100011000","010100000",8,'1'); -- (1, 2, 0, 2, 1, 1, 0, 0, 0)
sync_reset;
check_mem(2941,"100011000","010100001",2,'1'); -- (1, 2, 0, 2, 1, 1, 0, 0, 2)
sync_reset;
check_mem(2942,"100011010","010100001",2,'1'); -- (1, 2, 0, 2, 1, 1, 0, 1, 2)
sync_reset;
check_mem(2943,"100011000","010100010",2,'1'); -- (1, 2, 0, 2, 1, 1, 0, 2, 0)
sync_reset;
check_mem(2944,"100011100","010100001",2,'1'); -- (1, 2, 0, 2, 1, 1, 1, 0, 2)
sync_reset;
check_mem(2945,"100011100","010100010",2,'1'); -- (1, 2, 0, 2, 1, 1, 1, 2, 0)
sync_reset;
check_mem(2946,"100011100","010100011",2,'1'); -- (1, 2, 0, 2, 1, 1, 1, 2, 2)
sync_reset;
check_mem(2947,"100011000","010100100",8,'1'); -- (1, 2, 0, 2, 1, 1, 2, 0, 0)
sync_reset;
check_mem(2948,"100011010","010100100",8,'1'); -- (1, 2, 0, 2, 1, 1, 2, 1, 0)
sync_reset;
check_mem(2949,"100011010","010100101",2,'1'); -- (1, 2, 0, 2, 1, 1, 2, 1, 2)
sync_reset;
check_mem(2950,"100010010","010101000",2,'1'); -- (1, 2, 0, 2, 1, 2, 0, 1, 0)
sync_reset;
check_mem(2951,"100010100","010101000",2,'1'); -- (1, 2, 0, 2, 1, 2, 1, 0, 0)
sync_reset;
check_mem(2952,"100010110","010101000",2,'1'); -- (1, 2, 0, 2, 1, 2, 1, 1, 0)
sync_reset;
check_mem(2953,"100010110","010101001",2,'1'); -- (1, 2, 0, 2, 1, 2, 1, 1, 2)
sync_reset;
check_mem(2954,"100000011","010110000",5,'1'); -- (1, 2, 0, 2, 2, 0, 0, 1, 1)
sync_reset;
check_mem(2955,"100000101","010110000",7,'1'); -- (1, 2, 0, 2, 2, 0, 1, 0, 1)
sync_reset;
check_mem(2956,"100000110","010110000",8,'1'); -- (1, 2, 0, 2, 2, 0, 1, 1, 0)
sync_reset;
check_mem(2957,"100001001","010110000",2,'1'); -- (1, 2, 0, 2, 2, 1, 0, 0, 1)
sync_reset;
check_mem(2958,"100001010","010110000",8,'1'); -- (1, 2, 0, 2, 2, 1, 0, 1, 0)
sync_reset;
check_mem(2959,"100001011","010110000",2,'1'); -- (1, 2, 0, 2, 2, 1, 0, 1, 1)
sync_reset;
check_mem(2960,"100001100","010110000",7,'1'); -- (1, 2, 0, 2, 2, 1, 1, 0, 0)
sync_reset;
check_mem(2961,"100001101","010110000",7,'1'); -- (1, 2, 0, 2, 2, 1, 1, 0, 1)
sync_reset;
check_mem(2962,"100001110","010110000",8,'1'); -- (1, 2, 0, 2, 2, 1, 1, 1, 0)
sync_reset;
check_mem(2963,"100001110","010110001",2,'1'); -- (1, 2, 0, 2, 2, 1, 1, 1, 2)
sync_reset;
check_mem(2964,"100001011","010110100",2,'1'); -- (1, 2, 0, 2, 2, 1, 2, 1, 1)
sync_reset;
check_mem(2965,"101000000","010000000",4,'1'); -- (1, 2, 1, 0, 0, 0, 0, 0, 0)
sync_reset;
check_mem(2966,"101000000","010000001",6,'1'); -- (1, 2, 1, 0, 0, 0, 0, 0, 2)
sync_reset;
check_mem(2967,"101000010","010000001",3,'1'); -- (1, 2, 1, 0, 0, 0, 0, 1, 2)
sync_reset;
check_mem(2968,"101000000","010000010",4,'1'); -- (1, 2, 1, 0, 0, 0, 0, 2, 0)
sync_reset;
check_mem(2969,"101000001","010000010",4,'1'); -- (1, 2, 1, 0, 0, 0, 0, 2, 1)
sync_reset;
check_mem(2970,"101000100","010000001",3,'1'); -- (1, 2, 1, 0, 0, 0, 1, 0, 2)
sync_reset;
check_mem(2971,"101000100","010000010",4,'1'); -- (1, 2, 1, 0, 0, 0, 1, 2, 0)
sync_reset;
check_mem(2972,"101000100","010000011",3,'1'); -- (1, 2, 1, 0, 0, 0, 1, 2, 2)
sync_reset;
check_mem(2973,"101000000","010000100",8,'1'); -- (1, 2, 1, 0, 0, 0, 2, 0, 0)
sync_reset;
check_mem(2974,"101000001","010000100",3,'1'); -- (1, 2, 1, 0, 0, 0, 2, 0, 1)
sync_reset;
check_mem(2975,"101000010","010000100",4,'1'); -- (1, 2, 1, 0, 0, 0, 2, 1, 0)
sync_reset;
check_mem(2976,"101000010","010000101",3,'1'); -- (1, 2, 1, 0, 0, 0, 2, 1, 2)
sync_reset;
check_mem(2977,"101000001","010000110",4,'1'); -- (1, 2, 1, 0, 0, 0, 2, 2, 1)
sync_reset;
check_mem(2978,"101001000","010000001",7,'1'); -- (1, 2, 1, 0, 0, 1, 0, 0, 2)
sync_reset;
check_mem(2979,"101001000","010000010",4,'1'); -- (1, 2, 1, 0, 0, 1, 0, 2, 0)
sync_reset;
check_mem(2980,"101001000","010000011",3,'1'); -- (1, 2, 1, 0, 0, 1, 0, 2, 2)
sync_reset;
check_mem(2981,"101001100","010000011",4,'1'); -- (1, 2, 1, 0, 0, 1, 1, 2, 2)
sync_reset;
check_mem(2982,"101001000","010000100",8,'1'); -- (1, 2, 1, 0, 0, 1, 2, 0, 0)
sync_reset;
check_mem(2983,"101001000","010000101",7,'1'); -- (1, 2, 1, 0, 0, 1, 2, 0, 2)
sync_reset;
check_mem(2984,"101001010","010000101",3,'1'); -- (1, 2, 1, 0, 0, 1, 2, 1, 2)
sync_reset;
check_mem(2985,"101001000","010000110",8,'1'); -- (1, 2, 1, 0, 0, 1, 2, 2, 0)
sync_reset;
check_mem(2986,"101000000","010001000",4,'1'); -- (1, 2, 1, 0, 0, 2, 0, 0, 0)
sync_reset;
check_mem(2987,"101000001","010001000",4,'1'); -- (1, 2, 1, 0, 0, 2, 0, 0, 1)
sync_reset;
check_mem(2988,"101000010","010001000",4,'1'); -- (1, 2, 1, 0, 0, 2, 0, 1, 0)
sync_reset;
check_mem(2989,"101000010","010001001",6,'1'); -- (1, 2, 1, 0, 0, 2, 0, 1, 2)
sync_reset;
check_mem(2990,"101000001","010001010",4,'1'); -- (1, 2, 1, 0, 0, 2, 0, 2, 1)
sync_reset;
check_mem(2991,"101000100","010001000",3,'1'); -- (1, 2, 1, 0, 0, 2, 1, 0, 0)
sync_reset;
check_mem(2992,"101000100","010001001",3,'1'); -- (1, 2, 1, 0, 0, 2, 1, 0, 2)
sync_reset;
check_mem(2993,"101000110","010001001",3,'1'); -- (1, 2, 1, 0, 0, 2, 1, 1, 2)
sync_reset;
check_mem(2994,"101000100","010001010",3,'1'); -- (1, 2, 1, 0, 0, 2, 1, 2, 0)
sync_reset;
check_mem(2995,"101000101","010001010",4,'1'); -- (1, 2, 1, 0, 0, 2, 1, 2, 1)
sync_reset;
check_mem(2996,"101000001","010001100",4,'1'); -- (1, 2, 1, 0, 0, 2, 2, 0, 1)
sync_reset;
check_mem(2997,"101000010","010001100",3,'1'); -- (1, 2, 1, 0, 0, 2, 2, 1, 0)
sync_reset;
check_mem(2998,"101000011","010001100",4,'1'); -- (1, 2, 1, 0, 0, 2, 2, 1, 1)
sync_reset;
check_mem(2999,"101010000","010000001",6,'1'); -- (1, 2, 1, 0, 1, 0, 0, 0, 2)
sync_reset;
check_mem(3000,"101010000","010000010",3,'1'); -- (1, 2, 1, 0, 1, 0, 0, 2, 0)
sync_reset;
check_mem(3001,"101010000","010000011",6,'1'); -- (1, 2, 1, 0, 1, 0, 0, 2, 2)
sync_reset;
check_mem(3002,"101010000","010000100",8,'1'); -- (1, 2, 1, 0, 1, 0, 2, 0, 0)
sync_reset;
check_mem(3003,"101010000","010000101",7,'1'); -- (1, 2, 1, 0, 1, 0, 2, 0, 2)
sync_reset;
check_mem(3004,"101010010","010000101",3,'1'); -- (1, 2, 1, 0, 1, 0, 2, 1, 2)
sync_reset;
check_mem(3005,"101010000","010000110",8,'1'); -- (1, 2, 1, 0, 1, 0, 2, 2, 0)
sync_reset;
check_mem(3006,"101011000","010000011",6,'1'); -- (1, 2, 1, 0, 1, 1, 0, 2, 2)
sync_reset;
check_mem(3007,"101011000","010000101",7,'1'); -- (1, 2, 1, 0, 1, 1, 2, 0, 2)
sync_reset;
check_mem(3008,"101011000","010000110",8,'1'); -- (1, 2, 1, 0, 1, 1, 2, 2, 0)
sync_reset;
check_mem(3009,"101010000","010001000",3,'1'); -- (1, 2, 1, 0, 1, 2, 0, 0, 0)
sync_reset;
check_mem(3010,"101010000","010001001",6,'1'); -- (1, 2, 1, 0, 1, 2, 0, 0, 2)
sync_reset;
check_mem(3011,"101010010","010001001",6,'1'); -- (1, 2, 1, 0, 1, 2, 0, 1, 2)
sync_reset;
check_mem(3012,"101010000","010001010",3,'1'); -- (1, 2, 1, 0, 1, 2, 0, 2, 0)
sync_reset;
check_mem(3013,"101010000","010001100",8,'1'); -- (1, 2, 1, 0, 1, 2, 2, 0, 0)
sync_reset;
check_mem(3014,"101010010","010001100",8,'1'); -- (1, 2, 1, 0, 1, 2, 2, 1, 0)
sync_reset;
check_mem(3015,"101010010","010001101",3,'1'); -- (1, 2, 1, 0, 1, 2, 2, 1, 2)
sync_reset;
check_mem(3016,"101000000","010010000",7,'1'); -- (1, 2, 1, 0, 2, 0, 0, 0, 0)
sync_reset;
check_mem(3017,"101000001","010010000",5,'1'); -- (1, 2, 1, 0, 2, 0, 0, 0, 1)
sync_reset;
check_mem(3018,"101000010","010010000",3,'1'); -- (1, 2, 1, 0, 2, 0, 0, 1, 0)
sync_reset;
check_mem(3019,"101000010","010010001",3,'1'); -- (1, 2, 1, 0, 2, 0, 0, 1, 2)
sync_reset;
check_mem(3020,"101000100","010010000",3,'1'); -- (1, 2, 1, 0, 2, 0, 1, 0, 0)
sync_reset;
check_mem(3021,"101000100","010010001",3,'1'); -- (1, 2, 1, 0, 2, 0, 1, 0, 2)
sync_reset;
check_mem(3022,"101000110","010010001",3,'1'); -- (1, 2, 1, 0, 2, 0, 1, 1, 2)
sync_reset;
check_mem(3023,"101000001","010010100",5,'1'); -- (1, 2, 1, 0, 2, 0, 2, 0, 1)
sync_reset;
check_mem(3024,"101000010","010010100",3,'1'); -- (1, 2, 1, 0, 2, 0, 2, 1, 0)
sync_reset;
check_mem(3025,"101000011","010010100",5,'1'); -- (1, 2, 1, 0, 2, 0, 2, 1, 1)
sync_reset;
check_mem(3026,"101001000","010010000",7,'1'); -- (1, 2, 1, 0, 2, 1, 0, 0, 0)
sync_reset;
check_mem(3027,"101001000","010010001",7,'1'); -- (1, 2, 1, 0, 2, 1, 0, 0, 2)
sync_reset;
check_mem(3028,"101001010","010010001",3,'1'); -- (1, 2, 1, 0, 2, 1, 0, 1, 2)
sync_reset;
check_mem(3029,"101001100","010010001",7,'1'); -- (1, 2, 1, 0, 2, 1, 1, 0, 2)
sync_reset;
check_mem(3030,"101001000","010010100",8,'1'); -- (1, 2, 1, 0, 2, 1, 2, 0, 0)
sync_reset;
check_mem(3031,"101001010","010010100",8,'1'); -- (1, 2, 1, 0, 2, 1, 2, 1, 0)
sync_reset;
check_mem(3032,"101001010","010010101",3,'1'); -- (1, 2, 1, 0, 2, 1, 2, 1, 2)
sync_reset;
check_mem(3033,"101000001","010011000",3,'1'); -- (1, 2, 1, 0, 2, 2, 0, 0, 1)
sync_reset;
check_mem(3034,"101000010","010011000",3,'1'); -- (1, 2, 1, 0, 2, 2, 0, 1, 0)
sync_reset;
check_mem(3035,"101000011","010011000",3,'1'); -- (1, 2, 1, 0, 2, 2, 0, 1, 1)
sync_reset;
check_mem(3036,"101000100","010011000",3,'1'); -- (1, 2, 1, 0, 2, 2, 1, 0, 0)
sync_reset;
check_mem(3037,"101000101","010011000",3,'1'); -- (1, 2, 1, 0, 2, 2, 1, 0, 1)
sync_reset;
check_mem(3038,"101000110","010011000",3,'1'); -- (1, 2, 1, 0, 2, 2, 1, 1, 0)
sync_reset;
check_mem(3039,"101000110","010011001",3,'1'); -- (1, 2, 1, 0, 2, 2, 1, 1, 2)
sync_reset;
check_mem(3040,"101000011","010011100",3,'1'); -- (1, 2, 1, 0, 2, 2, 2, 1, 1)
sync_reset;
check_mem(3041,"101100000","010000001",6,'1'); -- (1, 2, 1, 1, 0, 0, 0, 0, 2)
sync_reset;
check_mem(3042,"101100000","010000010",4,'1'); -- (1, 2, 1, 1, 0, 0, 0, 2, 0)
sync_reset;
check_mem(3043,"101100000","010000011",6,'1'); -- (1, 2, 1, 1, 0, 0, 0, 2, 2)
sync_reset;
check_mem(3044,"101100000","010000100",7,'1'); -- (1, 2, 1, 1, 0, 0, 2, 0, 0)
sync_reset;
check_mem(3045,"101100000","010000101",7,'1'); -- (1, 2, 1, 1, 0, 0, 2, 0, 2)
sync_reset;
check_mem(3046,"101100010","010000101",4,'1'); -- (1, 2, 1, 1, 0, 0, 2, 1, 2)
sync_reset;
check_mem(3047,"101100000","010000110",4,'1'); -- (1, 2, 1, 1, 0, 0, 2, 2, 0)
sync_reset;
check_mem(3048,"101100001","010000110",4,'1'); -- (1, 2, 1, 1, 0, 0, 2, 2, 1)
sync_reset;
check_mem(3049,"101101000","010000011",4,'1'); -- (1, 2, 1, 1, 0, 1, 0, 2, 2)
sync_reset;
check_mem(3050,"101101000","010000101",7,'1'); -- (1, 2, 1, 1, 0, 1, 2, 0, 2)
sync_reset;
check_mem(3051,"101101000","010000110",4,'1'); -- (1, 2, 1, 1, 0, 1, 2, 2, 0)
sync_reset;
check_mem(3052,"101100000","010001000",6,'1'); -- (1, 2, 1, 1, 0, 2, 0, 0, 0)
sync_reset;
check_mem(3053,"101100000","010001001",6,'1'); -- (1, 2, 1, 1, 0, 2, 0, 0, 2)
sync_reset;
check_mem(3054,"101100010","010001001",6,'1'); -- (1, 2, 1, 1, 0, 2, 0, 1, 2)
sync_reset;
check_mem(3055,"101100000","010001010",4,'1'); -- (1, 2, 1, 1, 0, 2, 0, 2, 0)
sync_reset;
check_mem(3056,"101100001","010001010",4,'1'); -- (1, 2, 1, 1, 0, 2, 0, 2, 1)
sync_reset;
check_mem(3057,"101100000","010001100",4,'1'); -- (1, 2, 1, 1, 0, 2, 2, 0, 0)
sync_reset;
check_mem(3058,"101100001","010001100",4,'1'); -- (1, 2, 1, 1, 0, 2, 2, 0, 1)
sync_reset;
check_mem(3059,"101100010","010001100",4,'1'); -- (1, 2, 1, 1, 0, 2, 2, 1, 0)
sync_reset;
check_mem(3060,"101100010","010001101",4,'1'); -- (1, 2, 1, 1, 0, 2, 2, 1, 2)
sync_reset;
check_mem(3061,"101100001","010001110",4,'1'); -- (1, 2, 1, 1, 0, 2, 2, 2, 1)
sync_reset;
check_mem(3062,"101110000","010000011",6,'1'); -- (1, 2, 1, 1, 1, 0, 0, 2, 2)
sync_reset;
check_mem(3063,"101110000","010000101",7,'1'); -- (1, 2, 1, 1, 1, 0, 2, 0, 2)
sync_reset;
check_mem(3064,"101110000","010000110",8,'1'); -- (1, 2, 1, 1, 1, 0, 2, 2, 0)
sync_reset;
check_mem(3065,"101110000","010001001",6,'1'); -- (1, 2, 1, 1, 1, 2, 0, 0, 2)
sync_reset;
check_mem(3066,"101110000","010001010",6,'1'); -- (1, 2, 1, 1, 1, 2, 0, 2, 0)
sync_reset;
check_mem(3067,"101110000","010001011",6,'1'); -- (1, 2, 1, 1, 1, 2, 0, 2, 2)
sync_reset;
check_mem(3068,"101110000","010001100",8,'1'); -- (1, 2, 1, 1, 1, 2, 2, 0, 0)
sync_reset;
check_mem(3069,"101110000","010001101",7,'1'); -- (1, 2, 1, 1, 1, 2, 2, 0, 2)
sync_reset;
check_mem(3070,"101110000","010001110",8,'1'); -- (1, 2, 1, 1, 1, 2, 2, 2, 0)
sync_reset;
check_mem(3071,"101100000","010010000",7,'1'); -- (1, 2, 1, 1, 2, 0, 0, 0, 0)
sync_reset;
check_mem(3072,"101100000","010010001",6,'1'); -- (1, 2, 1, 1, 2, 0, 0, 0, 2)
sync_reset;
check_mem(3073,"101100010","010010001",6,'1'); -- (1, 2, 1, 1, 2, 0, 0, 1, 2)
sync_reset;
check_mem(3074,"101100000","010010100",7,'1'); -- (1, 2, 1, 1, 2, 0, 2, 0, 0)
sync_reset;
check_mem(3075,"101100001","010010100",7,'1'); -- (1, 2, 1, 1, 2, 0, 2, 0, 1)
sync_reset;
check_mem(3076,"101100010","010010100",5,'1'); -- (1, 2, 1, 1, 2, 0, 2, 1, 0)
sync_reset;
check_mem(3077,"101100010","010010101",5,'1'); -- (1, 2, 1, 1, 2, 0, 2, 1, 2)
sync_reset;
check_mem(3078,"101101000","010010001",7,'1'); -- (1, 2, 1, 1, 2, 1, 0, 0, 2)
sync_reset;
check_mem(3079,"101101000","010010100",7,'1'); -- (1, 2, 1, 1, 2, 1, 2, 0, 0)
sync_reset;
check_mem(3080,"101101000","010010101",7,'1'); -- (1, 2, 1, 1, 2, 1, 2, 0, 2)
sync_reset;
check_mem(3081,"101100000","010011000",6,'1'); -- (1, 2, 1, 1, 2, 2, 0, 0, 0)
sync_reset;
check_mem(3082,"101100001","010011000",7,'1'); -- (1, 2, 1, 1, 2, 2, 0, 0, 1)
sync_reset;
check_mem(3083,"101100010","010011000",6,'1'); -- (1, 2, 1, 1, 2, 2, 0, 1, 0)
sync_reset;
check_mem(3084,"101100010","010011001",6,'1'); -- (1, 2, 1, 1, 2, 2, 0, 1, 2)
sync_reset;
check_mem(3085,"101100001","010011100",7,'1'); -- (1, 2, 1, 1, 2, 2, 2, 0, 1)
sync_reset;
check_mem(3086,"101100010","010011100",8,'1'); -- (1, 2, 1, 1, 2, 2, 2, 1, 0)
sync_reset;
check_mem(3087,"101000000","010100000",4,'1'); -- (1, 2, 1, 2, 0, 0, 0, 0, 0)
sync_reset;
check_mem(3088,"101000001","010100000",4,'1'); -- (1, 2, 1, 2, 0, 0, 0, 0, 1)
sync_reset;
check_mem(3089,"101000010","010100000",4,'1'); -- (1, 2, 1, 2, 0, 0, 0, 1, 0)
sync_reset;
check_mem(3090,"101000010","010100001",4,'1'); -- (1, 2, 1, 2, 0, 0, 0, 1, 2)
sync_reset;
check_mem(3091,"101000001","010100010",4,'1'); -- (1, 2, 1, 2, 0, 0, 0, 2, 1)
sync_reset;
check_mem(3092,"101000100","010100000",4,'1'); -- (1, 2, 1, 2, 0, 0, 1, 0, 0)
sync_reset;
check_mem(3093,"101000100","010100001",4,'1'); -- (1, 2, 1, 2, 0, 0, 1, 0, 2)
sync_reset;
check_mem(3094,"101000110","010100001",4,'1'); -- (1, 2, 1, 2, 0, 0, 1, 1, 2)
sync_reset;
check_mem(3095,"101000100","010100010",4,'1'); -- (1, 2, 1, 2, 0, 0, 1, 2, 0)
sync_reset;
check_mem(3096,"101000101","010100010",4,'1'); -- (1, 2, 1, 2, 0, 0, 1, 2, 1)
sync_reset;
check_mem(3097,"101000001","010100100",4,'1'); -- (1, 2, 1, 2, 0, 0, 2, 0, 1)
sync_reset;
check_mem(3098,"101000010","010100100",8,'1'); -- (1, 2, 1, 2, 0, 0, 2, 1, 0)
sync_reset;
check_mem(3099,"101000011","010100100",4,'1'); -- (1, 2, 1, 2, 0, 0, 2, 1, 1)
sync_reset;
check_mem(3100,"101001000","010100000",8,'1'); -- (1, 2, 1, 2, 0, 1, 0, 0, 0)
sync_reset;
check_mem(3101,"101001000","010100001",4,'1'); -- (1, 2, 1, 2, 0, 1, 0, 0, 2)
sync_reset;
check_mem(3102,"101001010","010100001",4,'1'); -- (1, 2, 1, 2, 0, 1, 0, 1, 2)
sync_reset;
check_mem(3103,"101001000","010100010",4,'1'); -- (1, 2, 1, 2, 0, 1, 0, 2, 0)
sync_reset;
check_mem(3104,"101001100","010100001",4,'1'); -- (1, 2, 1, 2, 0, 1, 1, 0, 2)
sync_reset;
check_mem(3105,"101001100","010100010",4,'1'); -- (1, 2, 1, 2, 0, 1, 1, 2, 0)
sync_reset;
check_mem(3106,"101001100","010100011",4,'1'); -- (1, 2, 1, 2, 0, 1, 1, 2, 2)
sync_reset;
check_mem(3107,"101001000","010100100",8,'1'); -- (1, 2, 1, 2, 0, 1, 2, 0, 0)
sync_reset;
check_mem(3108,"101001010","010100100",8,'1'); -- (1, 2, 1, 2, 0, 1, 2, 1, 0)
sync_reset;
check_mem(3109,"101001010","010100101",4,'1'); -- (1, 2, 1, 2, 0, 1, 2, 1, 2)
sync_reset;
check_mem(3110,"101000001","010101000",4,'1'); -- (1, 2, 1, 2, 0, 2, 0, 0, 1)
sync_reset;
check_mem(3111,"101000010","010101000",4,'1'); -- (1, 2, 1, 2, 0, 2, 0, 1, 0)
sync_reset;
check_mem(3112,"101000011","010101000",4,'1'); -- (1, 2, 1, 2, 0, 2, 0, 1, 1)
sync_reset;
check_mem(3113,"101000100","010101000",4,'1'); -- (1, 2, 1, 2, 0, 2, 1, 0, 0)
sync_reset;
check_mem(3114,"101000101","010101000",4,'1'); -- (1, 2, 1, 2, 0, 2, 1, 0, 1)
sync_reset;
check_mem(3115,"101000110","010101000",4,'1'); -- (1, 2, 1, 2, 0, 2, 1, 1, 0)
sync_reset;
check_mem(3116,"101000110","010101001",4,'1'); -- (1, 2, 1, 2, 0, 2, 1, 1, 2)
sync_reset;
check_mem(3117,"101000101","010101010",4,'1'); -- (1, 2, 1, 2, 0, 2, 1, 2, 1)
sync_reset;
check_mem(3118,"101000011","010101100",4,'1'); -- (1, 2, 1, 2, 0, 2, 2, 1, 1)
sync_reset;
check_mem(3119,"101010000","010100000",5,'1'); -- (1, 2, 1, 2, 1, 0, 0, 0, 0)
sync_reset;
check_mem(3120,"101010000","010100001",6,'1'); -- (1, 2, 1, 2, 1, 0, 0, 0, 2)
sync_reset;
check_mem(3121,"101010010","010100001",6,'1'); -- (1, 2, 1, 2, 1, 0, 0, 1, 2)
sync_reset;
check_mem(3122,"101010000","010100010",5,'1'); -- (1, 2, 1, 2, 1, 0, 0, 2, 0)
sync_reset;
check_mem(3123,"101010000","010100100",8,'1'); -- (1, 2, 1, 2, 1, 0, 2, 0, 0)
sync_reset;
check_mem(3124,"101010010","010100100",8,'1'); -- (1, 2, 1, 2, 1, 0, 2, 1, 0)
sync_reset;
check_mem(3125,"101010010","010100101",5,'1'); -- (1, 2, 1, 2, 1, 0, 2, 1, 2)
sync_reset;
check_mem(3126,"101011000","010100001",6,'1'); -- (1, 2, 1, 2, 1, 1, 0, 0, 2)
sync_reset;
check_mem(3127,"101011000","010100010",6,'1'); -- (1, 2, 1, 2, 1, 1, 0, 2, 0)
sync_reset;
check_mem(3128,"101011000","010100011",6,'1'); -- (1, 2, 1, 2, 1, 1, 0, 2, 2)
sync_reset;
check_mem(3129,"101011000","010100100",8,'1'); -- (1, 2, 1, 2, 1, 1, 2, 0, 0)
sync_reset;
check_mem(3130,"101011000","010100101",7,'1'); -- (1, 2, 1, 2, 1, 1, 2, 0, 2)
sync_reset;
check_mem(3131,"101011000","010100110",8,'1'); -- (1, 2, 1, 2, 1, 1, 2, 2, 0)
sync_reset;
check_mem(3132,"101010000","010101000",6,'1'); -- (1, 2, 1, 2, 1, 2, 0, 0, 0)
sync_reset;
check_mem(3133,"101010010","010101000",6,'1'); -- (1, 2, 1, 2, 1, 2, 0, 1, 0)
sync_reset;
check_mem(3134,"101010010","010101001",6,'1'); -- (1, 2, 1, 2, 1, 2, 0, 1, 2)
sync_reset;
check_mem(3135,"101010010","010101100",8,'1'); -- (1, 2, 1, 2, 1, 2, 2, 1, 0)
sync_reset;
check_mem(3136,"101000001","010110000",5,'1'); -- (1, 2, 1, 2, 2, 0, 0, 0, 1)
sync_reset;
check_mem(3137,"101000010","010110000",5,'1'); -- (1, 2, 1, 2, 2, 0, 0, 1, 0)
sync_reset;
check_mem(3138,"101000011","010110000",5,'1'); -- (1, 2, 1, 2, 2, 0, 0, 1, 1)
sync_reset;
check_mem(3139,"101000100","010110000",5,'1'); -- (1, 2, 1, 2, 2, 0, 1, 0, 0)
sync_reset;
check_mem(3140,"101000101","010110000",5,'1'); -- (1, 2, 1, 2, 2, 0, 1, 0, 1)
sync_reset;
check_mem(3141,"101000110","010110000",5,'1'); -- (1, 2, 1, 2, 2, 0, 1, 1, 0)
sync_reset;
check_mem(3142,"101000110","010110001",5,'1'); -- (1, 2, 1, 2, 2, 0, 1, 1, 2)
sync_reset;
check_mem(3143,"101000011","010110100",5,'1'); -- (1, 2, 1, 2, 2, 0, 2, 1, 1)
sync_reset;
check_mem(3144,"101001000","010110000",8,'1'); -- (1, 2, 1, 2, 2, 1, 0, 0, 0)
sync_reset;
check_mem(3145,"101001010","010110000",8,'1'); -- (1, 2, 1, 2, 2, 1, 0, 1, 0)
sync_reset;
check_mem(3146,"101001010","010110001",6,'1'); -- (1, 2, 1, 2, 2, 1, 0, 1, 2)
sync_reset;
check_mem(3147,"101001100","010110000",7,'1'); -- (1, 2, 1, 2, 2, 1, 1, 0, 0)
sync_reset;
check_mem(3148,"101001100","010110001",7,'1'); -- (1, 2, 1, 2, 2, 1, 1, 0, 2)
sync_reset;
check_mem(3149,"101001010","010110100",8,'1'); -- (1, 2, 1, 2, 2, 1, 2, 1, 0)
sync_reset;
check_mem(3150,"100000001","011000000",3,'1'); -- (1, 2, 2, 0, 0, 0, 0, 0, 1)
sync_reset;
check_mem(3151,"100000010","011000000",3,'1'); -- (1, 2, 2, 0, 0, 0, 0, 1, 0)
sync_reset;
check_mem(3152,"100000011","011000000",3,'1'); -- (1, 2, 2, 0, 0, 0, 0, 1, 1)
sync_reset;
check_mem(3153,"100000100","011000000",3,'1'); -- (1, 2, 2, 0, 0, 0, 1, 0, 0)
sync_reset;
check_mem(3154,"100000101","011000000",3,'1'); -- (1, 2, 2, 0, 0, 0, 1, 0, 1)
sync_reset;
check_mem(3155,"100000110","011000000",3,'1'); -- (1, 2, 2, 0, 0, 0, 1, 1, 0)
sync_reset;
check_mem(3156,"100000110","011000001",3,'1'); -- (1, 2, 2, 0, 0, 0, 1, 1, 2)
sync_reset;
check_mem(3157,"100000101","011000010",3,'1'); -- (1, 2, 2, 0, 0, 0, 1, 2, 1)
sync_reset;
check_mem(3158,"100000011","011000100",4,'1'); -- (1, 2, 2, 0, 0, 0, 2, 1, 1)
sync_reset;
check_mem(3159,"100001000","011000000",3,'1'); -- (1, 2, 2, 0, 0, 1, 0, 0, 0)
sync_reset;
check_mem(3160,"100001001","011000000",4,'1'); -- (1, 2, 2, 0, 0, 1, 0, 0, 1)
sync_reset;
check_mem(3161,"100001010","011000000",3,'1'); -- (1, 2, 2, 0, 0, 1, 0, 1, 0)
sync_reset;
check_mem(3162,"100001010","011000001",3,'1'); -- (1, 2, 2, 0, 0, 1, 0, 1, 2)
sync_reset;
check_mem(3163,"100001001","011000010",4,'1'); -- (1, 2, 2, 0, 0, 1, 0, 2, 1)
sync_reset;
check_mem(3164,"100001100","011000000",3,'1'); -- (1, 2, 2, 0, 0, 1, 1, 0, 0)
sync_reset;
check_mem(3165,"100001100","011000001",3,'1'); -- (1, 2, 2, 0, 0, 1, 1, 0, 2)
sync_reset;
check_mem(3166,"100001110","011000001",3,'1'); -- (1, 2, 2, 0, 0, 1, 1, 1, 2)
sync_reset;
check_mem(3167,"100001100","011000010",3,'1'); -- (1, 2, 2, 0, 0, 1, 1, 2, 0)
sync_reset;
check_mem(3168,"100001101","011000010",4,'1'); -- (1, 2, 2, 0, 0, 1, 1, 2, 1)
sync_reset;
check_mem(3169,"100001001","011000100",4,'1'); -- (1, 2, 2, 0, 0, 1, 2, 0, 1)
sync_reset;
check_mem(3170,"100001010","011000100",4,'1'); -- (1, 2, 2, 0, 0, 1, 2, 1, 0)
sync_reset;
check_mem(3171,"100001011","011000100",4,'1'); -- (1, 2, 2, 0, 0, 1, 2, 1, 1)
sync_reset;
check_mem(3172,"100000011","011001000",3,'1'); -- (1, 2, 2, 0, 0, 2, 0, 1, 1)
sync_reset;
check_mem(3173,"100000101","011001000",3,'1'); -- (1, 2, 2, 0, 0, 2, 1, 0, 1)
sync_reset;
check_mem(3174,"100000110","011001000",3,'1'); -- (1, 2, 2, 0, 0, 2, 1, 1, 0)
sync_reset;
check_mem(3175,"100010000","011000000",3,'1'); -- (1, 2, 2, 0, 1, 0, 0, 0, 0)
sync_reset;
check_mem(3176,"100010010","011000000",8,'1'); -- (1, 2, 2, 0, 1, 0, 0, 1, 0)
sync_reset;
check_mem(3177,"100010010","011000001",5,'1'); -- (1, 2, 2, 0, 1, 0, 0, 1, 2)
sync_reset;
check_mem(3178,"100010100","011000000",3,'1'); -- (1, 2, 2, 0, 1, 0, 1, 0, 0)
sync_reset;
check_mem(3179,"100010100","011000001",3,'1'); -- (1, 2, 2, 0, 1, 0, 1, 0, 2)
sync_reset;
check_mem(3180,"100010110","011000001",5,'1'); -- (1, 2, 2, 0, 1, 0, 1, 1, 2)
sync_reset;
check_mem(3181,"100010100","011000010",3,'1'); -- (1, 2, 2, 0, 1, 0, 1, 2, 0)
sync_reset;
check_mem(3182,"100010010","011000100",3,'1'); -- (1, 2, 2, 0, 1, 0, 2, 1, 0)
sync_reset;
check_mem(3183,"100011000","011000000",3,'1'); -- (1, 2, 2, 0, 1, 1, 0, 0, 0)
sync_reset;
check_mem(3184,"100011000","011000001",3,'1'); -- (1, 2, 2, 0, 1, 1, 0, 0, 2)
sync_reset;
check_mem(3185,"100011010","011000001",3,'1'); -- (1, 2, 2, 0, 1, 1, 0, 1, 2)
sync_reset;
check_mem(3186,"100011000","011000010",3,'1'); -- (1, 2, 2, 0, 1, 1, 0, 2, 0)
sync_reset;
check_mem(3187,"100011100","011000001",3,'1'); -- (1, 2, 2, 0, 1, 1, 1, 0, 2)
sync_reset;
check_mem(3188,"100011100","011000010",3,'1'); -- (1, 2, 2, 0, 1, 1, 1, 2, 0)
sync_reset;
check_mem(3189,"100011100","011000011",3,'1'); -- (1, 2, 2, 0, 1, 1, 1, 2, 2)
sync_reset;
check_mem(3190,"100011000","011000100",3,'1'); -- (1, 2, 2, 0, 1, 1, 2, 0, 0)
sync_reset;
check_mem(3191,"100011010","011000100",3,'1'); -- (1, 2, 2, 0, 1, 1, 2, 1, 0)
sync_reset;
check_mem(3192,"100011010","011000101",3,'1'); -- (1, 2, 2, 0, 1, 1, 2, 1, 2)
sync_reset;
check_mem(3193,"100010010","011001000",8,'1'); -- (1, 2, 2, 0, 1, 2, 0, 1, 0)
sync_reset;
check_mem(3194,"100010100","011001000",3,'1'); -- (1, 2, 2, 0, 1, 2, 1, 0, 0)
sync_reset;
check_mem(3195,"100010110","011001000",8,'1'); -- (1, 2, 2, 0, 1, 2, 1, 1, 0)
sync_reset;
check_mem(3196,"100000011","011010000",6,'1'); -- (1, 2, 2, 0, 2, 0, 0, 1, 1)
sync_reset;
check_mem(3197,"100000101","011010000",3,'1'); -- (1, 2, 2, 0, 2, 0, 1, 0, 1)
sync_reset;
check_mem(3198,"100000110","011010000",3,'1'); -- (1, 2, 2, 0, 2, 0, 1, 1, 0)
sync_reset;
check_mem(3199,"100001001","011010000",3,'1'); -- (1, 2, 2, 0, 2, 1, 0, 0, 1)
sync_reset;
check_mem(3200,"100001010","011010000",6,'1'); -- (1, 2, 2, 0, 2, 1, 0, 1, 0)
sync_reset;
check_mem(3201,"100001011","011010000",6,'1'); -- (1, 2, 2, 0, 2, 1, 0, 1, 1)
sync_reset;
check_mem(3202,"100001100","011010000",3,'1'); -- (1, 2, 2, 0, 2, 1, 1, 0, 0)
sync_reset;
check_mem(3203,"100001101","011010000",7,'1'); -- (1, 2, 2, 0, 2, 1, 1, 0, 1)
sync_reset;
check_mem(3204,"100001110","011010000",3,'1'); -- (1, 2, 2, 0, 2, 1, 1, 1, 0)
sync_reset;
check_mem(3205,"100001110","011010001",3,'1'); -- (1, 2, 2, 0, 2, 1, 1, 1, 2)
sync_reset;
check_mem(3206,"100100000","011000000",4,'1'); -- (1, 2, 2, 1, 0, 0, 0, 0, 0)
sync_reset;
check_mem(3207,"100100001","011000000",4,'1'); -- (1, 2, 2, 1, 0, 0, 0, 0, 1)
sync_reset;
check_mem(3208,"100100010","011000000",4,'1'); -- (1, 2, 2, 1, 0, 0, 0, 1, 0)
sync_reset;
check_mem(3209,"100100010","011000001",5,'1'); -- (1, 2, 2, 1, 0, 0, 0, 1, 2)
sync_reset;
check_mem(3210,"100100001","011000010",4,'1'); -- (1, 2, 2, 1, 0, 0, 0, 2, 1)
sync_reset;
check_mem(3211,"100100001","011000100",4,'1'); -- (1, 2, 2, 1, 0, 0, 2, 0, 1)
sync_reset;
check_mem(3212,"100100010","011000100",4,'1'); -- (1, 2, 2, 1, 0, 0, 2, 1, 0)
sync_reset;
check_mem(3213,"100100011","011000100",4,'1'); -- (1, 2, 2, 1, 0, 0, 2, 1, 1)
sync_reset;
check_mem(3214,"100101000","011000000",4,'1'); -- (1, 2, 2, 1, 0, 1, 0, 0, 0)
sync_reset;
check_mem(3215,"100101000","011000001",4,'1'); -- (1, 2, 2, 1, 0, 1, 0, 0, 2)
sync_reset;
check_mem(3216,"100101010","011000001",4,'1'); -- (1, 2, 2, 1, 0, 1, 0, 1, 2)
sync_reset;
check_mem(3217,"100101000","011000010",4,'1'); -- (1, 2, 2, 1, 0, 1, 0, 2, 0)
sync_reset;
check_mem(3218,"100101001","011000010",4,'1'); -- (1, 2, 2, 1, 0, 1, 0, 2, 1)
sync_reset;
check_mem(3219,"100101000","011000100",4,'1'); -- (1, 2, 2, 1, 0, 1, 2, 0, 0)
sync_reset;
check_mem(3220,"100101001","011000100",4,'1'); -- (1, 2, 2, 1, 0, 1, 2, 0, 1)
sync_reset;
check_mem(3221,"100101010","011000100",4,'1'); -- (1, 2, 2, 1, 0, 1, 2, 1, 0)
sync_reset;
check_mem(3222,"100101010","011000101",4,'1'); -- (1, 2, 2, 1, 0, 1, 2, 1, 2)
sync_reset;
check_mem(3223,"100101001","011000110",4,'1'); -- (1, 2, 2, 1, 0, 1, 2, 2, 1)
sync_reset;
check_mem(3224,"100100001","011001000",4,'1'); -- (1, 2, 2, 1, 0, 2, 0, 0, 1)
sync_reset;
check_mem(3225,"100100010","011001000",6,'1'); -- (1, 2, 2, 1, 0, 2, 0, 1, 0)
sync_reset;
check_mem(3226,"100100011","011001000",4,'1'); -- (1, 2, 2, 1, 0, 2, 0, 1, 1)
sync_reset;
check_mem(3227,"100100011","011001100",4,'1'); -- (1, 2, 2, 1, 0, 2, 2, 1, 1)
sync_reset;
check_mem(3228,"100110000","011000000",5,'1'); -- (1, 2, 2, 1, 1, 0, 0, 0, 0)
sync_reset;
check_mem(3229,"100110000","011000001",5,'1'); -- (1, 2, 2, 1, 1, 0, 0, 0, 2)
sync_reset;
check_mem(3230,"100110010","011000001",5,'1'); -- (1, 2, 2, 1, 1, 0, 0, 1, 2)
sync_reset;
check_mem(3231,"100110000","011000010",5,'1'); -- (1, 2, 2, 1, 1, 0, 0, 2, 0)
sync_reset;
check_mem(3232,"100110000","011000100",5,'1'); -- (1, 2, 2, 1, 1, 0, 2, 0, 0)
sync_reset;
check_mem(3233,"100110010","011000100",5,'1'); -- (1, 2, 2, 1, 1, 0, 2, 1, 0)
sync_reset;
check_mem(3234,"100110010","011000101",5,'1'); -- (1, 2, 2, 1, 1, 0, 2, 1, 2)
sync_reset;
check_mem(3235,"100110000","011001000",6,'1'); -- (1, 2, 2, 1, 1, 2, 0, 0, 0)
sync_reset;
check_mem(3236,"100110010","011001000",8,'1'); -- (1, 2, 2, 1, 1, 2, 0, 1, 0)
sync_reset;
check_mem(3237,"100110010","011001100",8,'1'); -- (1, 2, 2, 1, 1, 2, 2, 1, 0)
sync_reset;
check_mem(3238,"100100001","011010000",6,'1'); -- (1, 2, 2, 1, 2, 0, 0, 0, 1)
sync_reset;
check_mem(3239,"100100010","011010000",6,'1'); -- (1, 2, 2, 1, 2, 0, 0, 1, 0)
sync_reset;
check_mem(3240,"100100011","011010000",6,'1'); -- (1, 2, 2, 1, 2, 0, 0, 1, 1)
sync_reset;
check_mem(3241,"100101000","011010000",6,'1'); -- (1, 2, 2, 1, 2, 1, 0, 0, 0)
sync_reset;
check_mem(3242,"100101001","011010000",6,'1'); -- (1, 2, 2, 1, 2, 1, 0, 0, 1)
sync_reset;
check_mem(3243,"100101010","011010000",6,'1'); -- (1, 2, 2, 1, 2, 1, 0, 1, 0)
sync_reset;
check_mem(3244,"100101010","011010001",6,'1'); -- (1, 2, 2, 1, 2, 1, 0, 1, 2)
sync_reset;
check_mem(3245,"100100011","011011000",6,'1'); -- (1, 2, 2, 1, 2, 2, 0, 1, 1)
sync_reset;
check_mem(3246,"100000011","011100000",4,'1'); -- (1, 2, 2, 2, 0, 0, 0, 1, 1)
sync_reset;
check_mem(3247,"100000101","011100000",4,'1'); -- (1, 2, 2, 2, 0, 0, 1, 0, 1)
sync_reset;
check_mem(3248,"100000110","011100000",8,'1'); -- (1, 2, 2, 2, 0, 0, 1, 1, 0)
sync_reset;
check_mem(3249,"100001001","011100000",4,'1'); -- (1, 2, 2, 2, 0, 1, 0, 0, 1)
sync_reset;
check_mem(3250,"100001010","011100000",8,'1'); -- (1, 2, 2, 2, 0, 1, 0, 1, 0)
sync_reset;
check_mem(3251,"100001011","011100000",4,'1'); -- (1, 2, 2, 2, 0, 1, 0, 1, 1)
sync_reset;
check_mem(3252,"100001100","011100000",8,'1'); -- (1, 2, 2, 2, 0, 1, 1, 0, 0)
sync_reset;
check_mem(3253,"100001101","011100000",4,'1'); -- (1, 2, 2, 2, 0, 1, 1, 0, 1)
sync_reset;
check_mem(3254,"100001110","011100000",8,'1'); -- (1, 2, 2, 2, 0, 1, 1, 1, 0)
sync_reset;
check_mem(3255,"100001110","011100001",4,'1'); -- (1, 2, 2, 2, 0, 1, 1, 1, 2)
sync_reset;
check_mem(3256,"100001101","011100010",4,'1'); -- (1, 2, 2, 2, 0, 1, 1, 2, 1)
sync_reset;
check_mem(3257,"100001011","011100100",4,'1'); -- (1, 2, 2, 2, 0, 1, 2, 1, 1)
sync_reset;
check_mem(3258,"100010010","011100000",8,'1'); -- (1, 2, 2, 2, 1, 0, 0, 1, 0)
sync_reset;
check_mem(3259,"100010100","011100000",8,'1'); -- (1, 2, 2, 2, 1, 0, 1, 0, 0)
sync_reset;
check_mem(3260,"100010110","011100000",8,'1'); -- (1, 2, 2, 2, 1, 0, 1, 1, 0)
sync_reset;
check_mem(3261,"100010110","011100001",5,'1'); -- (1, 2, 2, 2, 1, 0, 1, 1, 2)
sync_reset;
check_mem(3262,"100011000","011100000",8,'1'); -- (1, 2, 2, 2, 1, 1, 0, 0, 0)
sync_reset;
check_mem(3263,"100011010","011100000",8,'1'); -- (1, 2, 2, 2, 1, 1, 0, 1, 0)
sync_reset;
check_mem(3264,"100011010","011100001",6,'1'); -- (1, 2, 2, 2, 1, 1, 0, 1, 2)
sync_reset;
check_mem(3265,"100011100","011100000",8,'1'); -- (1, 2, 2, 2, 1, 1, 1, 0, 0)
sync_reset;
check_mem(3266,"100011100","011100001",7,'1'); -- (1, 2, 2, 2, 1, 1, 1, 0, 2)
sync_reset;
check_mem(3267,"100011100","011100010",8,'1'); -- (1, 2, 2, 2, 1, 1, 1, 2, 0)
sync_reset;
check_mem(3268,"100011010","011100100",8,'1'); -- (1, 2, 2, 2, 1, 1, 2, 1, 0)
sync_reset;
check_mem(3269,"100010110","011101000",8,'1'); -- (1, 2, 2, 2, 1, 2, 1, 1, 0)
sync_reset;
check_mem(3270,"100001011","011110000",6,'1'); -- (1, 2, 2, 2, 2, 1, 0, 1, 1)
sync_reset;
check_mem(3271,"100001101","011110000",7,'1'); -- (1, 2, 2, 2, 2, 1, 1, 0, 1)
sync_reset;
check_mem(3272,"100001110","011110000",8,'1'); -- (1, 2, 2, 2, 2, 1, 1, 1, 0)
sync_reset;
check_mem(3273,"000000001","100000000",2,'1'); -- (2, 0, 0, 0, 0, 0, 0, 0, 1)
sync_reset;
check_mem(3274,"000000010","100000000",6,'1'); -- (2, 0, 0, 0, 0, 0, 0, 1, 0)
sync_reset;
check_mem(3275,"000000011","100000000",6,'1'); -- (2, 0, 0, 0, 0, 0, 0, 1, 1)
sync_reset;
check_mem(3276,"000000100","100000000",2,'1'); -- (2, 0, 0, 0, 0, 0, 1, 0, 0)
sync_reset;
check_mem(3277,"000000101","100000000",1,'1'); -- (2, 0, 0, 0, 0, 0, 1, 0, 1)
sync_reset;
check_mem(3278,"000000110","100000000",1,'1'); -- (2, 0, 0, 0, 0, 0, 1, 1, 0)
sync_reset;
check_mem(3279,"000000110","100000001",4,'1'); -- (2, 0, 0, 0, 0, 0, 1, 1, 2)
sync_reset;
check_mem(3280,"000000101","100000010",2,'1'); -- (2, 0, 0, 0, 0, 0, 1, 2, 1)
sync_reset;
check_mem(3281,"000000011","100000100",1,'1'); -- (2, 0, 0, 0, 0, 0, 2, 1, 1)
sync_reset;
check_mem(3282,"000001000","100000000",2,'1'); -- (2, 0, 0, 0, 0, 1, 0, 0, 0)
sync_reset;
check_mem(3283,"000001001","100000000",2,'1'); -- (2, 0, 0, 0, 0, 1, 0, 0, 1)
sync_reset;
check_mem(3284,"000001010","100000000",2,'1'); -- (2, 0, 0, 0, 0, 1, 0, 1, 0)
sync_reset;
check_mem(3285,"000001010","100000001",4,'1'); -- (2, 0, 0, 0, 0, 1, 0, 1, 2)
sync_reset;
check_mem(3286,"000001001","100000010",2,'1'); -- (2, 0, 0, 0, 0, 1, 0, 2, 1)
sync_reset;
check_mem(3287,"000001100","100000000",2,'1'); -- (2, 0, 0, 0, 0, 1, 1, 0, 0)
sync_reset;
check_mem(3288,"000001100","100000001",4,'1'); -- (2, 0, 0, 0, 0, 1, 1, 0, 2)
sync_reset;
check_mem(3289,"000001110","100000001",1,'1'); -- (2, 0, 0, 0, 0, 1, 1, 1, 2)
sync_reset;
check_mem(3290,"000001100","100000010",2,'1'); -- (2, 0, 0, 0, 0, 1, 1, 2, 0)
sync_reset;
check_mem(3291,"000001101","100000010",2,'1'); -- (2, 0, 0, 0, 0, 1, 1, 2, 1)
sync_reset;
check_mem(3292,"000001001","100000100",2,'1'); -- (2, 0, 0, 0, 0, 1, 2, 0, 1)
sync_reset;
check_mem(3293,"000001010","100000100",1,'1'); -- (2, 0, 0, 0, 0, 1, 2, 1, 0)
sync_reset;
check_mem(3294,"000001011","100000100",2,'1'); -- (2, 0, 0, 0, 0, 1, 2, 1, 1)
sync_reset;
check_mem(3295,"000000011","100001000",1,'1'); -- (2, 0, 0, 0, 0, 2, 0, 1, 1)
sync_reset;
check_mem(3296,"000000101","100001000",2,'1'); -- (2, 0, 0, 0, 0, 2, 1, 0, 1)
sync_reset;
check_mem(3297,"000000110","100001000",1,'1'); -- (2, 0, 0, 0, 0, 2, 1, 1, 0)
sync_reset;
check_mem(3298,"000010000","100000000",1,'1'); -- (2, 0, 0, 0, 1, 0, 0, 0, 0)
sync_reset;
check_mem(3299,"000010001","100000000",2,'1'); -- (2, 0, 0, 0, 1, 0, 0, 0, 1)
sync_reset;
check_mem(3300,"000010010","100000000",1,'1'); -- (2, 0, 0, 0, 1, 0, 0, 1, 0)
sync_reset;
check_mem(3301,"000010010","100000001",1,'1'); -- (2, 0, 0, 0, 1, 0, 0, 1, 2)
sync_reset;
check_mem(3302,"000010001","100000010",2,'1'); -- (2, 0, 0, 0, 1, 0, 0, 2, 1)
sync_reset;
check_mem(3303,"000010100","100000000",2,'1'); -- (2, 0, 0, 0, 1, 0, 1, 0, 0)
sync_reset;
check_mem(3304,"000010100","100000001",1,'1'); -- (2, 0, 0, 0, 1, 0, 1, 0, 2)
sync_reset;
check_mem(3305,"000010110","100000001",1,'1'); -- (2, 0, 0, 0, 1, 0, 1, 1, 2)
sync_reset;
check_mem(3306,"000010100","100000010",2,'1'); -- (2, 0, 0, 0, 1, 0, 1, 2, 0)
sync_reset;
check_mem(3307,"000010101","100000010",2,'1'); -- (2, 0, 0, 0, 1, 0, 1, 2, 1)
sync_reset;
check_mem(3308,"000010001","100000100",3,'1'); -- (2, 0, 0, 0, 1, 0, 2, 0, 1)
sync_reset;
check_mem(3309,"000010010","100000100",1,'1'); -- (2, 0, 0, 0, 1, 0, 2, 1, 0)
sync_reset;
check_mem(3310,"000010011","100000100",1,'1'); -- (2, 0, 0, 0, 1, 0, 2, 1, 1)
sync_reset;
check_mem(3311,"000011000","100000000",3,'1'); -- (2, 0, 0, 0, 1, 1, 0, 0, 0)
sync_reset;
check_mem(3312,"000011000","100000001",1,'1'); -- (2, 0, 0, 0, 1, 1, 0, 0, 2)
sync_reset;
check_mem(3313,"000011010","100000001",1,'1'); -- (2, 0, 0, 0, 1, 1, 0, 1, 2)
sync_reset;
check_mem(3314,"000011000","100000010",2,'1'); -- (2, 0, 0, 0, 1, 1, 0, 2, 0)
sync_reset;
check_mem(3315,"000011001","100000010",1,'1'); -- (2, 0, 0, 0, 1, 1, 0, 2, 1)
sync_reset;
check_mem(3316,"000011100","100000001",1,'1'); -- (2, 0, 0, 0, 1, 1, 1, 0, 2)
sync_reset;
check_mem(3317,"000011100","100000010",1,'1'); -- (2, 0, 0, 0, 1, 1, 1, 2, 0)
sync_reset;
check_mem(3318,"000011100","100000011",1,'1'); -- (2, 0, 0, 0, 1, 1, 1, 2, 2)
sync_reset;
check_mem(3319,"000011000","100000100",3,'1'); -- (2, 0, 0, 0, 1, 1, 2, 0, 0)
sync_reset;
check_mem(3320,"000011001","100000100",3,'1'); -- (2, 0, 0, 0, 1, 1, 2, 0, 1)
sync_reset;
check_mem(3321,"000011010","100000100",3,'1'); -- (2, 0, 0, 0, 1, 1, 2, 1, 0)
sync_reset;
check_mem(3322,"000011010","100000101",1,'1'); -- (2, 0, 0, 0, 1, 1, 2, 1, 2)
sync_reset;
check_mem(3323,"000011001","100000110",2,'1'); -- (2, 0, 0, 0, 1, 1, 2, 2, 1)
sync_reset;
check_mem(3324,"000010001","100001000",6,'1'); -- (2, 0, 0, 0, 1, 2, 0, 0, 1)
sync_reset;
check_mem(3325,"000010010","100001000",1,'1'); -- (2, 0, 0, 0, 1, 2, 0, 1, 0)
sync_reset;
check_mem(3326,"000010011","100001000",1,'1'); -- (2, 0, 0, 0, 1, 2, 0, 1, 1)
sync_reset;
check_mem(3327,"000010100","100001000",1,'1'); -- (2, 0, 0, 0, 1, 2, 1, 0, 0)
sync_reset;
check_mem(3328,"000010101","100001000",1,'1'); -- (2, 0, 0, 0, 1, 2, 1, 0, 1)
sync_reset;
check_mem(3329,"000010110","100001000",1,'1'); -- (2, 0, 0, 0, 1, 2, 1, 1, 0)
sync_reset;
check_mem(3330,"000010110","100001001",1,'1'); -- (2, 0, 0, 0, 1, 2, 1, 1, 2)
sync_reset;
check_mem(3331,"000010101","100001010",2,'1'); -- (2, 0, 0, 0, 1, 2, 1, 2, 1)
sync_reset;
check_mem(3332,"000010011","100001100",1,'1'); -- (2, 0, 0, 0, 1, 2, 2, 1, 1)
sync_reset;
check_mem(3333,"000000011","100010000",2,'1'); -- (2, 0, 0, 0, 2, 0, 0, 1, 1)
sync_reset;
check_mem(3334,"000000101","100010000",2,'1'); -- (2, 0, 0, 0, 2, 0, 1, 0, 1)
sync_reset;
check_mem(3335,"000000110","100010000",8,'1'); -- (2, 0, 0, 0, 2, 0, 1, 1, 0)
sync_reset;
check_mem(3336,"000001001","100010000",2,'1'); -- (2, 0, 0, 0, 2, 1, 0, 0, 1)
sync_reset;
check_mem(3337,"000001010","100010000",8,'1'); -- (2, 0, 0, 0, 2, 1, 0, 1, 0)
sync_reset;
check_mem(3338,"000001011","100010000",1,'1'); -- (2, 0, 0, 0, 2, 1, 0, 1, 1)
sync_reset;
check_mem(3339,"000001100","100010000",8,'1'); -- (2, 0, 0, 0, 2, 1, 1, 0, 0)
sync_reset;
check_mem(3340,"000001101","100010000",1,'1'); -- (2, 0, 0, 0, 2, 1, 1, 0, 1)
sync_reset;
check_mem(3341,"000001110","100010000",8,'1'); -- (2, 0, 0, 0, 2, 1, 1, 1, 0)
sync_reset;
check_mem(3342,"000001101","100010010",2,'1'); -- (2, 0, 0, 0, 2, 1, 1, 2, 1)
sync_reset;
check_mem(3343,"000001011","100010100",2,'1'); -- (2, 0, 0, 0, 2, 1, 2, 1, 1)
sync_reset;
check_mem(3344,"000100000","100000000",1,'1'); -- (2, 0, 0, 1, 0, 0, 0, 0, 0)
sync_reset;
check_mem(3345,"000100001","100000000",2,'1'); -- (2, 0, 0, 1, 0, 0, 0, 0, 1)
sync_reset;
check_mem(3346,"000100010","100000000",2,'1'); -- (2, 0, 0, 1, 0, 0, 0, 1, 0)
sync_reset;
check_mem(3347,"000100010","100000001",4,'1'); -- (2, 0, 0, 1, 0, 0, 0, 1, 2)
sync_reset;
check_mem(3348,"000100001","100000010",5,'1'); -- (2, 0, 0, 1, 0, 0, 0, 2, 1)
sync_reset;
check_mem(3349,"000100100","100000000",1,'1'); -- (2, 0, 0, 1, 0, 0, 1, 0, 0)
sync_reset;
check_mem(3350,"000100100","100000001",4,'1'); -- (2, 0, 0, 1, 0, 0, 1, 0, 2)
sync_reset;
check_mem(3351,"000100110","100000001",1,'1'); -- (2, 0, 0, 1, 0, 0, 1, 1, 2)
sync_reset;
check_mem(3352,"000100100","100000010",4,'1'); -- (2, 0, 0, 1, 0, 0, 1, 2, 0)
sync_reset;
check_mem(3353,"000100101","100000010",1,'1'); -- (2, 0, 0, 1, 0, 0, 1, 2, 1)
sync_reset;
check_mem(3354,"000100001","100000100",5,'1'); -- (2, 0, 0, 1, 0, 0, 2, 0, 1)
sync_reset;
check_mem(3355,"000100010","100000100",4,'1'); -- (2, 0, 0, 1, 0, 0, 2, 1, 0)
sync_reset;
check_mem(3356,"000100011","100000100",2,'1'); -- (2, 0, 0, 1, 0, 0, 2, 1, 1)
sync_reset;
check_mem(3357,"000101000","100000000",4,'1'); -- (2, 0, 0, 1, 0, 1, 0, 0, 0)
sync_reset;
check_mem(3358,"000101000","100000001",4,'1'); -- (2, 0, 0, 1, 0, 1, 0, 0, 2)
sync_reset;
check_mem(3359,"000101010","100000001",4,'1'); -- (2, 0, 0, 1, 0, 1, 0, 1, 2)
sync_reset;
check_mem(3360,"000101000","100000010",2,'1'); -- (2, 0, 0, 1, 0, 1, 0, 2, 0)
sync_reset;
check_mem(3361,"000101001","100000010",1,'1'); -- (2, 0, 0, 1, 0, 1, 0, 2, 1)
sync_reset;
check_mem(3362,"000101100","100000001",4,'1'); -- (2, 0, 0, 1, 0, 1, 1, 0, 2)
sync_reset;
check_mem(3363,"000101100","100000010",4,'1'); -- (2, 0, 0, 1, 0, 1, 1, 2, 0)
sync_reset;
check_mem(3364,"000101100","100000011",4,'1'); -- (2, 0, 0, 1, 0, 1, 1, 2, 2)
sync_reset;
check_mem(3365,"000101000","100000100",2,'1'); -- (2, 0, 0, 1, 0, 1, 2, 0, 0)
sync_reset;
check_mem(3366,"000101001","100000100",1,'1'); -- (2, 0, 0, 1, 0, 1, 2, 0, 1)
sync_reset;
check_mem(3367,"000101010","100000100",4,'1'); -- (2, 0, 0, 1, 0, 1, 2, 1, 0)
sync_reset;
check_mem(3368,"000101010","100000101",4,'1'); -- (2, 0, 0, 1, 0, 1, 2, 1, 2)
sync_reset;
check_mem(3369,"000101001","100000110",1,'1'); -- (2, 0, 0, 1, 0, 1, 2, 2, 1)
sync_reset;
check_mem(3370,"000100001","100001000",1,'1'); -- (2, 0, 0, 1, 0, 2, 0, 0, 1)
sync_reset;
check_mem(3371,"000100010","100001000",1,'1'); -- (2, 0, 0, 1, 0, 2, 0, 1, 0)
sync_reset;
check_mem(3372,"000100011","100001000",6,'1'); -- (2, 0, 0, 1, 0, 2, 0, 1, 1)
sync_reset;
check_mem(3373,"000100100","100001000",2,'1'); -- (2, 0, 0, 1, 0, 2, 1, 0, 0)
sync_reset;
check_mem(3374,"000100101","100001000",7,'1'); -- (2, 0, 0, 1, 0, 2, 1, 0, 1)
sync_reset;
check_mem(3375,"000100110","100001000",8,'1'); -- (2, 0, 0, 1, 0, 2, 1, 1, 0)
sync_reset;
check_mem(3376,"000100110","100001001",1,'1'); -- (2, 0, 0, 1, 0, 2, 1, 1, 2)
sync_reset;
check_mem(3377,"000100101","100001010",1,'1'); -- (2, 0, 0, 1, 0, 2, 1, 2, 1)
sync_reset;
check_mem(3378,"000100011","100001100",1,'1'); -- (2, 0, 0, 1, 0, 2, 2, 1, 1)
sync_reset;
check_mem(3379,"000110000","100000000",5,'1'); -- (2, 0, 0, 1, 1, 0, 0, 0, 0)
sync_reset;
check_mem(3380,"000110000","100000001",1,'1'); -- (2, 0, 0, 1, 1, 0, 0, 0, 2)
sync_reset;
check_mem(3381,"000110010","100000001",1,'1'); -- (2, 0, 0, 1, 1, 0, 0, 1, 2)
sync_reset;
check_mem(3382,"000110000","100000010",2,'1'); -- (2, 0, 0, 1, 1, 0, 0, 2, 0)
sync_reset;
check_mem(3383,"000110001","100000010",5,'1'); -- (2, 0, 0, 1, 1, 0, 0, 2, 1)
sync_reset;
check_mem(3384,"000110100","100000001",1,'1'); -- (2, 0, 0, 1, 1, 0, 1, 0, 2)
sync_reset;
check_mem(3385,"000110100","100000010",1,'1'); -- (2, 0, 0, 1, 1, 0, 1, 2, 0)
sync_reset;
check_mem(3386,"000110100","100000011",1,'1'); -- (2, 0, 0, 1, 1, 0, 1, 2, 2)
sync_reset;
check_mem(3387,"000110000","100000100",1,'1'); -- (2, 0, 0, 1, 1, 0, 2, 0, 0)
sync_reset;
check_mem(3388,"000110001","100000100",5,'1'); -- (2, 0, 0, 1, 1, 0, 2, 0, 1)
sync_reset;
check_mem(3389,"000110010","100000100",1,'1'); -- (2, 0, 0, 1, 1, 0, 2, 1, 0)
sync_reset;
check_mem(3390,"000110010","100000101",1,'1'); -- (2, 0, 0, 1, 1, 0, 2, 1, 2)
sync_reset;
check_mem(3391,"000110001","100000110",5,'1'); -- (2, 0, 0, 1, 1, 0, 2, 2, 1)
sync_reset;
check_mem(3392,"000110000","100001000",1,'1'); -- (2, 0, 0, 1, 1, 2, 0, 0, 0)
sync_reset;
check_mem(3393,"000110001","100001000",1,'1'); -- (2, 0, 0, 1, 1, 2, 0, 0, 1)
sync_reset;
check_mem(3394,"000110010","100001000",1,'1'); -- (2, 0, 0, 1, 1, 2, 0, 1, 0)
sync_reset;
check_mem(3395,"000110010","100001001",1,'1'); -- (2, 0, 0, 1, 1, 2, 0, 1, 2)
sync_reset;
check_mem(3396,"000110001","100001010",1,'1'); -- (2, 0, 0, 1, 1, 2, 0, 2, 1)
sync_reset;
check_mem(3397,"000110100","100001000",2,'1'); -- (2, 0, 0, 1, 1, 2, 1, 0, 0)
sync_reset;
check_mem(3398,"000110100","100001001",2,'1'); -- (2, 0, 0, 1, 1, 2, 1, 0, 2)
sync_reset;
check_mem(3399,"000110110","100001001",2,'1'); -- (2, 0, 0, 1, 1, 2, 1, 1, 2)
sync_reset;
check_mem(3400,"000110100","100001010",2,'1'); -- (2, 0, 0, 1, 1, 2, 1, 2, 0)
sync_reset;
check_mem(3401,"000110101","100001010",2,'1'); -- (2, 0, 0, 1, 1, 2, 1, 2, 1)
sync_reset;
check_mem(3402,"000110001","100001100",1,'1'); -- (2, 0, 0, 1, 1, 2, 2, 0, 1)
sync_reset;
check_mem(3403,"000110010","100001100",1,'1'); -- (2, 0, 0, 1, 1, 2, 2, 1, 0)
sync_reset;
check_mem(3404,"000110011","100001100",1,'1'); -- (2, 0, 0, 1, 1, 2, 2, 1, 1)
sync_reset;
check_mem(3405,"000100001","100010000",1,'1'); -- (2, 0, 0, 1, 2, 0, 0, 0, 1)
sync_reset;
check_mem(3406,"000100010","100010000",8,'1'); -- (2, 0, 0, 1, 2, 0, 0, 1, 0)
sync_reset;
check_mem(3407,"000100011","100010000",6,'1'); -- (2, 0, 0, 1, 2, 0, 0, 1, 1)
sync_reset;
check_mem(3408,"000100100","100010000",8,'1'); -- (2, 0, 0, 1, 2, 0, 1, 0, 0)
sync_reset;
check_mem(3409,"000100101","100010000",7,'1'); -- (2, 0, 0, 1, 2, 0, 1, 0, 1)
sync_reset;
check_mem(3410,"000100110","100010000",8,'1'); -- (2, 0, 0, 1, 2, 0, 1, 1, 0)
sync_reset;
check_mem(3411,"000100101","100010010",1,'1'); -- (2, 0, 0, 1, 2, 0, 1, 2, 1)
sync_reset;
check_mem(3412,"000100011","100010100",2,'1'); -- (2, 0, 0, 1, 2, 0, 2, 1, 1)
sync_reset;
check_mem(3413,"000101000","100010000",1,'1'); -- (2, 0, 0, 1, 2, 1, 0, 0, 0)
sync_reset;
check_mem(3414,"000101001","100010000",2,'1'); -- (2, 0, 0, 1, 2, 1, 0, 0, 1)
sync_reset;
check_mem(3415,"000101010","100010000",1,'1'); -- (2, 0, 0, 1, 2, 1, 0, 1, 0)
sync_reset;
check_mem(3416,"000101001","100010010",2,'1'); -- (2, 0, 0, 1, 2, 1, 0, 2, 1)
sync_reset;
check_mem(3417,"000101100","100010000",1,'1'); -- (2, 0, 0, 1, 2, 1, 1, 0, 0)
sync_reset;
check_mem(3418,"000101100","100010010",1,'1'); -- (2, 0, 0, 1, 2, 1, 1, 2, 0)
sync_reset;
check_mem(3419,"000101101","100010010",1,'1'); -- (2, 0, 0, 1, 2, 1, 1, 2, 1)
sync_reset;
check_mem(3420,"000101001","100010100",2,'1'); -- (2, 0, 0, 1, 2, 1, 2, 0, 1)
sync_reset;
check_mem(3421,"000101010","100010100",1,'1'); -- (2, 0, 0, 1, 2, 1, 2, 1, 0)
sync_reset;
check_mem(3422,"000101011","100010100",2,'1'); -- (2, 0, 0, 1, 2, 1, 2, 1, 1)
sync_reset;
check_mem(3423,"000100011","100011000",6,'1'); -- (2, 0, 0, 1, 2, 2, 0, 1, 1)
sync_reset;
check_mem(3424,"000100101","100011000",7,'1'); -- (2, 0, 0, 1, 2, 2, 1, 0, 1)
sync_reset;
check_mem(3425,"000100110","100011000",8,'1'); -- (2, 0, 0, 1, 2, 2, 1, 1, 0)
sync_reset;
check_mem(3426,"000000011","100100000",6,'1'); -- (2, 0, 0, 2, 0, 0, 0, 1, 1)
sync_reset;
check_mem(3427,"000000101","100100000",1,'1'); -- (2, 0, 0, 2, 0, 0, 1, 0, 1)
sync_reset;
check_mem(3428,"000000110","100100000",1,'1'); -- (2, 0, 0, 2, 0, 0, 1, 1, 0)
sync_reset;
check_mem(3429,"000001001","100100000",2,'1'); -- (2, 0, 0, 2, 0, 1, 0, 0, 1)
sync_reset;
check_mem(3430,"000001010","100100000",6,'1'); -- (2, 0, 0, 2, 0, 1, 0, 1, 0)
sync_reset;
check_mem(3431,"000001011","100100000",6,'1'); -- (2, 0, 0, 2, 0, 1, 0, 1, 1)
sync_reset;
check_mem(3432,"000001100","100100000",1,'1'); -- (2, 0, 0, 2, 0, 1, 1, 0, 0)
sync_reset;
check_mem(3433,"000001101","100100000",1,'1'); -- (2, 0, 0, 2, 0, 1, 1, 0, 1)
sync_reset;
check_mem(3434,"000001110","100100000",1,'1'); -- (2, 0, 0, 2, 0, 1, 1, 1, 0)
sync_reset;
check_mem(3435,"000001110","100100001",4,'1'); -- (2, 0, 0, 2, 0, 1, 1, 1, 2)
sync_reset;
check_mem(3436,"000001101","100100010",2,'1'); -- (2, 0, 0, 2, 0, 1, 1, 2, 1)
sync_reset;
check_mem(3437,"000010001","100100000",6,'1'); -- (2, 0, 0, 2, 1, 0, 0, 0, 1)
sync_reset;
check_mem(3438,"000010010","100100000",1,'1'); -- (2, 0, 0, 2, 1, 0, 0, 1, 0)
sync_reset;
check_mem(3439,"000010011","100100000",6,'1'); -- (2, 0, 0, 2, 1, 0, 0, 1, 1)
sync_reset;
check_mem(3440,"000010100","100100000",1,'1'); -- (2, 0, 0, 2, 1, 0, 1, 0, 0)
sync_reset;
check_mem(3441,"000010101","100100000",1,'1'); -- (2, 0, 0, 2, 1, 0, 1, 0, 1)
sync_reset;
check_mem(3442,"000010110","100100000",1,'1'); -- (2, 0, 0, 2, 1, 0, 1, 1, 0)
sync_reset;
check_mem(3443,"000010110","100100001",1,'1'); -- (2, 0, 0, 2, 1, 0, 1, 1, 2)
sync_reset;
check_mem(3444,"000010101","100100010",2,'1'); -- (2, 0, 0, 2, 1, 0, 1, 2, 1)
sync_reset;
check_mem(3445,"000011000","100100000",6,'1'); -- (2, 0, 0, 2, 1, 1, 0, 0, 0)
sync_reset;
check_mem(3446,"000011001","100100000",2,'1'); -- (2, 0, 0, 2, 1, 1, 0, 0, 1)
sync_reset;
check_mem(3447,"000011010","100100000",1,'1'); -- (2, 0, 0, 2, 1, 1, 0, 1, 0)
sync_reset;
check_mem(3448,"000011010","100100001",1,'1'); -- (2, 0, 0, 2, 1, 1, 0, 1, 2)
sync_reset;
check_mem(3449,"000011001","100100010",2,'1'); -- (2, 0, 0, 2, 1, 1, 0, 2, 1)
sync_reset;
check_mem(3450,"000011100","100100000",2,'1'); -- (2, 0, 0, 2, 1, 1, 1, 0, 0)
sync_reset;
check_mem(3451,"000011100","100100001",1,'1'); -- (2, 0, 0, 2, 1, 1, 1, 0, 2)
sync_reset;
check_mem(3452,"000011110","100100001",1,'1'); -- (2, 0, 0, 2, 1, 1, 1, 1, 2)
sync_reset;
check_mem(3453,"000011100","100100010",2,'1'); -- (2, 0, 0, 2, 1, 1, 1, 2, 0)
sync_reset;
check_mem(3454,"000011101","100100010",2,'1'); -- (2, 0, 0, 2, 1, 1, 1, 2, 1)
sync_reset;
check_mem(3455,"000010011","100101000",1,'1'); -- (2, 0, 0, 2, 1, 2, 0, 1, 1)
sync_reset;
check_mem(3456,"000010101","100101000",1,'1'); -- (2, 0, 0, 2, 1, 2, 1, 0, 1)
sync_reset;
check_mem(3457,"000010110","100101000",1,'1'); -- (2, 0, 0, 2, 1, 2, 1, 1, 0)
sync_reset;
check_mem(3458,"000001011","100110000",2,'1'); -- (2, 0, 0, 2, 2, 1, 0, 1, 1)
sync_reset;
check_mem(3459,"000001101","100110000",1,'1'); -- (2, 0, 0, 2, 2, 1, 1, 0, 1)
sync_reset;
check_mem(3460,"000001110","100110000",8,'1'); -- (2, 0, 0, 2, 2, 1, 1, 1, 0)
sync_reset;
check_mem(3461,"001000000","100000000",5,'1'); -- (2, 0, 1, 0, 0, 0, 0, 0, 0)
sync_reset;
check_mem(3462,"001000001","100000000",1,'1'); -- (2, 0, 1, 0, 0, 0, 0, 0, 1)
sync_reset;
check_mem(3463,"001000010","100000000",6,'1'); -- (2, 0, 1, 0, 0, 0, 0, 1, 0)
sync_reset;
check_mem(3464,"001000010","100000001",4,'1'); -- (2, 0, 1, 0, 0, 0, 0, 1, 2)
sync_reset;
check_mem(3465,"001000001","100000010",4,'1'); -- (2, 0, 1, 0, 0, 0, 0, 2, 1)
sync_reset;
check_mem(3466,"001000100","100000000",1,'1'); -- (2, 0, 1, 0, 0, 0, 1, 0, 0)
sync_reset;
check_mem(3467,"001000100","100000001",4,'1'); -- (2, 0, 1, 0, 0, 0, 1, 0, 2)
sync_reset;
check_mem(3468,"001000110","100000001",4,'1'); -- (2, 0, 1, 0, 0, 0, 1, 1, 2)
sync_reset;
check_mem(3469,"001000100","100000010",4,'1'); -- (2, 0, 1, 0, 0, 0, 1, 2, 0)
sync_reset;
check_mem(3470,"001000101","100000010",1,'1'); -- (2, 0, 1, 0, 0, 0, 1, 2, 1)
sync_reset;
check_mem(3471,"001000001","100000100",5,'1'); -- (2, 0, 1, 0, 0, 0, 2, 0, 1)
sync_reset;
check_mem(3472,"001000010","100000100",3,'1'); -- (2, 0, 1, 0, 0, 0, 2, 1, 0)
sync_reset;
check_mem(3473,"001000011","100000100",3,'1'); -- (2, 0, 1, 0, 0, 0, 2, 1, 1)
sync_reset;
check_mem(3474,"001001000","100000000",1,'1'); -- (2, 0, 1, 0, 0, 1, 0, 0, 0)
sync_reset;
check_mem(3475,"001001000","100000001",4,'1'); -- (2, 0, 1, 0, 0, 1, 0, 0, 2)
sync_reset;
check_mem(3476,"001001010","100000001",3,'1'); -- (2, 0, 1, 0, 0, 1, 0, 1, 2)
sync_reset;
check_mem(3477,"001001000","100000010",3,'1'); -- (2, 0, 1, 0, 0, 1, 0, 2, 0)
sync_reset;
check_mem(3478,"001001100","100000001",4,'1'); -- (2, 0, 1, 0, 0, 1, 1, 0, 2)
sync_reset;
check_mem(3479,"001001100","100000010",1,'1'); -- (2, 0, 1, 0, 0, 1, 1, 2, 0)
sync_reset;
check_mem(3480,"001001100","100000011",4,'1'); -- (2, 0, 1, 0, 0, 1, 1, 2, 2)
sync_reset;
check_mem(3481,"001001000","100000100",3,'1'); -- (2, 0, 1, 0, 0, 1, 2, 0, 0)
sync_reset;
check_mem(3482,"001001010","100000100",3,'1'); -- (2, 0, 1, 0, 0, 1, 2, 1, 0)
sync_reset;
check_mem(3483,"001001010","100000101",1,'1'); -- (2, 0, 1, 0, 0, 1, 2, 1, 2)
sync_reset;
check_mem(3484,"001000001","100001000",6,'1'); -- (2, 0, 1, 0, 0, 2, 0, 0, 1)
sync_reset;
check_mem(3485,"001000010","100001000",4,'1'); -- (2, 0, 1, 0, 0, 2, 0, 1, 0)
sync_reset;
check_mem(3486,"001000011","100001000",6,'1'); -- (2, 0, 1, 0, 0, 2, 0, 1, 1)
sync_reset;
check_mem(3487,"001000100","100001000",4,'1'); -- (2, 0, 1, 0, 0, 2, 1, 0, 0)
sync_reset;
check_mem(3488,"001000101","100001000",1,'1'); -- (2, 0, 1, 0, 0, 2, 1, 0, 1)
sync_reset;
check_mem(3489,"001000110","100001000",1,'1'); -- (2, 0, 1, 0, 0, 2, 1, 1, 0)
sync_reset;
check_mem(3490,"001000110","100001001",4,'1'); -- (2, 0, 1, 0, 0, 2, 1, 1, 2)
sync_reset;
check_mem(3491,"001000101","100001010",4,'1'); -- (2, 0, 1, 0, 0, 2, 1, 2, 1)
sync_reset;
check_mem(3492,"001000011","100001100",3,'1'); -- (2, 0, 1, 0, 0, 2, 2, 1, 1)
sync_reset;
check_mem(3493,"001010000","100000000",6,'1'); -- (2, 0, 1, 0, 1, 0, 0, 0, 0)
sync_reset;
check_mem(3494,"001010000","100000001",1,'1'); -- (2, 0, 1, 0, 1, 0, 0, 0, 2)
sync_reset;
check_mem(3495,"001010010","100000001",1,'1'); -- (2, 0, 1, 0, 1, 0, 0, 1, 2)
sync_reset;
check_mem(3496,"001010000","100000010",3,'1'); -- (2, 0, 1, 0, 1, 0, 0, 2, 0)
sync_reset;
check_mem(3497,"001010001","100000010",1,'1'); -- (2, 0, 1, 0, 1, 0, 0, 2, 1)
sync_reset;
check_mem(3498,"001010000","100000100",3,'1'); -- (2, 0, 1, 0, 1, 0, 2, 0, 0)
sync_reset;
check_mem(3499,"001010001","100000100",3,'1'); -- (2, 0, 1, 0, 1, 0, 2, 0, 1)
sync_reset;
check_mem(3500,"001010010","100000100",3,'1'); -- (2, 0, 1, 0, 1, 0, 2, 1, 0)
sync_reset;
check_mem(3501,"001010010","100000101",1,'1'); -- (2, 0, 1, 0, 1, 0, 2, 1, 2)
sync_reset;
check_mem(3502,"001010001","100000110",5,'1'); -- (2, 0, 1, 0, 1, 0, 2, 2, 1)
sync_reset;
check_mem(3503,"001011000","100000001",1,'1'); -- (2, 0, 1, 0, 1, 1, 0, 0, 2)
sync_reset;
check_mem(3504,"001011000","100000010",1,'1'); -- (2, 0, 1, 0, 1, 1, 0, 2, 0)
sync_reset;
check_mem(3505,"001011000","100000011",3,'1'); -- (2, 0, 1, 0, 1, 1, 0, 2, 2)
sync_reset;
check_mem(3506,"001011000","100000100",3,'1'); -- (2, 0, 1, 0, 1, 1, 2, 0, 0)
sync_reset;
check_mem(3507,"001011000","100000101",3,'1'); -- (2, 0, 1, 0, 1, 1, 2, 0, 2)
sync_reset;
check_mem(3508,"001011010","100000101",3,'1'); -- (2, 0, 1, 0, 1, 1, 2, 1, 2)
sync_reset;
check_mem(3509,"001011000","100000110",3,'1'); -- (2, 0, 1, 0, 1, 1, 2, 2, 0)
sync_reset;
check_mem(3510,"001010000","100001000",1,'1'); -- (2, 0, 1, 0, 1, 2, 0, 0, 0)
sync_reset;
check_mem(3511,"001010001","100001000",6,'1'); -- (2, 0, 1, 0, 1, 2, 0, 0, 1)
sync_reset;
check_mem(3512,"001010010","100001000",1,'1'); -- (2, 0, 1, 0, 1, 2, 0, 1, 0)
sync_reset;
check_mem(3513,"001010010","100001001",1,'1'); -- (2, 0, 1, 0, 1, 2, 0, 1, 2)
sync_reset;
check_mem(3514,"001010001","100001010",6,'1'); -- (2, 0, 1, 0, 1, 2, 0, 2, 1)
sync_reset;
check_mem(3515,"001010001","100001100",3,'1'); -- (2, 0, 1, 0, 1, 2, 2, 0, 1)
sync_reset;
check_mem(3516,"001010010","100001100",1,'1'); -- (2, 0, 1, 0, 1, 2, 2, 1, 0)
sync_reset;
check_mem(3517,"001010011","100001100",3,'1'); -- (2, 0, 1, 0, 1, 2, 2, 1, 1)
sync_reset;
check_mem(3518,"001000001","100010000",5,'1'); -- (2, 0, 1, 0, 2, 0, 0, 0, 1)
sync_reset;
check_mem(3519,"001000010","100010000",8,'1'); -- (2, 0, 1, 0, 2, 0, 0, 1, 0)
sync_reset;
check_mem(3520,"001000011","100010000",1,'1'); -- (2, 0, 1, 0, 2, 0, 0, 1, 1)
sync_reset;
check_mem(3521,"001000100","100010000",8,'1'); -- (2, 0, 1, 0, 2, 0, 1, 0, 0)
sync_reset;
check_mem(3522,"001000101","100010000",1,'1'); -- (2, 0, 1, 0, 2, 0, 1, 0, 1)
sync_reset;
check_mem(3523,"001000110","100010000",8,'1'); -- (2, 0, 1, 0, 2, 0, 1, 1, 0)
sync_reset;
check_mem(3524,"001000101","100010010",5,'1'); -- (2, 0, 1, 0, 2, 0, 1, 2, 1)
sync_reset;
check_mem(3525,"001000011","100010100",5,'1'); -- (2, 0, 1, 0, 2, 0, 2, 1, 1)
sync_reset;
check_mem(3526,"001001000","100010000",8,'1'); -- (2, 0, 1, 0, 2, 1, 0, 0, 0)
sync_reset;
check_mem(3527,"001001010","100010000",8,'1'); -- (2, 0, 1, 0, 2, 1, 0, 1, 0)
sync_reset;
check_mem(3528,"001001100","100010000",8,'1'); -- (2, 0, 1, 0, 2, 1, 1, 0, 0)
sync_reset;
check_mem(3529,"001001100","100010010",8,'1'); -- (2, 0, 1, 0, 2, 1, 1, 2, 0)
sync_reset;
check_mem(3530,"001001010","100010100",8,'1'); -- (2, 0, 1, 0, 2, 1, 2, 1, 0)
sync_reset;
check_mem(3531,"001000011","100011000",6,'1'); -- (2, 0, 1, 0, 2, 2, 0, 1, 1)
sync_reset;
check_mem(3532,"001000101","100011000",7,'1'); -- (2, 0, 1, 0, 2, 2, 1, 0, 1)
sync_reset;
check_mem(3533,"001000110","100011000",8,'1'); -- (2, 0, 1, 0, 2, 2, 1, 1, 0)
sync_reset;
check_mem(3534,"001100000","100000000",4,'1'); -- (2, 0, 1, 1, 0, 0, 0, 0, 0)
sync_reset;
check_mem(3535,"001100000","100000001",4,'1'); -- (2, 0, 1, 1, 0, 0, 0, 0, 2)
sync_reset;
check_mem(3536,"001100010","100000001",4,'1'); -- (2, 0, 1, 1, 0, 0, 0, 1, 2)
sync_reset;
check_mem(3537,"001100000","100000010",4,'1'); -- (2, 0, 1, 1, 0, 0, 0, 2, 0)
sync_reset;
check_mem(3538,"001100001","100000010",5,'1'); -- (2, 0, 1, 1, 0, 0, 0, 2, 1)
sync_reset;
check_mem(3539,"001100100","100000001",4,'1'); -- (2, 0, 1, 1, 0, 0, 1, 0, 2)
sync_reset;
check_mem(3540,"001100100","100000010",4,'1'); -- (2, 0, 1, 1, 0, 0, 1, 2, 0)
sync_reset;
check_mem(3541,"001100100","100000011",4,'1'); -- (2, 0, 1, 1, 0, 0, 1, 2, 2)
sync_reset;
check_mem(3542,"001100000","100000100",5,'1'); -- (2, 0, 1, 1, 0, 0, 2, 0, 0)
sync_reset;
check_mem(3543,"001100001","100000100",5,'1'); -- (2, 0, 1, 1, 0, 0, 2, 0, 1)
sync_reset;
check_mem(3544,"001100010","100000100",4,'1'); -- (2, 0, 1, 1, 0, 0, 2, 1, 0)
sync_reset;
check_mem(3545,"001100010","100000101",4,'1'); -- (2, 0, 1, 1, 0, 0, 2, 1, 2)
sync_reset;
check_mem(3546,"001100001","100000110",5,'1'); -- (2, 0, 1, 1, 0, 0, 2, 2, 1)
sync_reset;
check_mem(3547,"001101000","100000001",4,'1'); -- (2, 0, 1, 1, 0, 1, 0, 0, 2)
sync_reset;
check_mem(3548,"001101000","100000010",1,'1'); -- (2, 0, 1, 1, 0, 1, 0, 2, 0)
sync_reset;
check_mem(3549,"001101000","100000011",4,'1'); -- (2, 0, 1, 1, 0, 1, 0, 2, 2)
sync_reset;
check_mem(3550,"001101100","100000011",4,'1'); -- (2, 0, 1, 1, 0, 1, 1, 2, 2)
sync_reset;
check_mem(3551,"001101000","100000100",1,'1'); -- (2, 0, 1, 1, 0, 1, 2, 0, 0)
sync_reset;
check_mem(3552,"001101000","100000101",4,'1'); -- (2, 0, 1, 1, 0, 1, 2, 0, 2)
sync_reset;
check_mem(3553,"001101010","100000101",4,'1'); -- (2, 0, 1, 1, 0, 1, 2, 1, 2)
sync_reset;
check_mem(3554,"001101000","100000110",4,'1'); -- (2, 0, 1, 1, 0, 1, 2, 2, 0)
sync_reset;
check_mem(3555,"001100000","100001000",1,'1'); -- (2, 0, 1, 1, 0, 2, 0, 0, 0)
sync_reset;
check_mem(3556,"001100001","100001000",4,'1'); -- (2, 0, 1, 1, 0, 2, 0, 0, 1)
sync_reset;
check_mem(3557,"001100010","100001000",4,'1'); -- (2, 0, 1, 1, 0, 2, 0, 1, 0)
sync_reset;
check_mem(3558,"001100010","100001001",4,'1'); -- (2, 0, 1, 1, 0, 2, 0, 1, 2)
sync_reset;
check_mem(3559,"001100001","100001010",1,'1'); -- (2, 0, 1, 1, 0, 2, 0, 2, 1)
sync_reset;
check_mem(3560,"001100100","100001000",4,'1'); -- (2, 0, 1, 1, 0, 2, 1, 0, 0)
sync_reset;
check_mem(3561,"001100100","100001001",4,'1'); -- (2, 0, 1, 1, 0, 2, 1, 0, 2)
sync_reset;
check_mem(3562,"001100110","100001001",4,'1'); -- (2, 0, 1, 1, 0, 2, 1, 1, 2)
sync_reset;
check_mem(3563,"001100100","100001010",4,'1'); -- (2, 0, 1, 1, 0, 2, 1, 2, 0)
sync_reset;
check_mem(3564,"001100101","100001010",4,'1'); -- (2, 0, 1, 1, 0, 2, 1, 2, 1)
sync_reset;
check_mem(3565,"001100001","100001100",1,'1'); -- (2, 0, 1, 1, 0, 2, 2, 0, 1)
sync_reset;
check_mem(3566,"001100010","100001100",1,'1'); -- (2, 0, 1, 1, 0, 2, 2, 1, 0)
sync_reset;
check_mem(3567,"001100011","100001100",1,'1'); -- (2, 0, 1, 1, 0, 2, 2, 1, 1)
sync_reset;
check_mem(3568,"001110000","100000001",1,'1'); -- (2, 0, 1, 1, 1, 0, 0, 0, 2)
sync_reset;
check_mem(3569,"001110000","100000010",1,'1'); -- (2, 0, 1, 1, 1, 0, 0, 2, 0)
sync_reset;
check_mem(3570,"001110000","100000011",5,'1'); -- (2, 0, 1, 1, 1, 0, 0, 2, 2)
sync_reset;
check_mem(3571,"001110000","100000100",5,'1'); -- (2, 0, 1, 1, 1, 0, 2, 0, 0)
sync_reset;
check_mem(3572,"001110000","100000101",5,'1'); -- (2, 0, 1, 1, 1, 0, 2, 0, 2)
sync_reset;
check_mem(3573,"001110010","100000101",1,'1'); -- (2, 0, 1, 1, 1, 0, 2, 1, 2)
sync_reset;
check_mem(3574,"001110000","100000110",5,'1'); -- (2, 0, 1, 1, 1, 0, 2, 2, 0)
sync_reset;
check_mem(3575,"001110001","100000110",5,'1'); -- (2, 0, 1, 1, 1, 0, 2, 2, 1)
sync_reset;
check_mem(3576,"001110000","100001000",6,'1'); -- (2, 0, 1, 1, 1, 2, 0, 0, 0)
sync_reset;
check_mem(3577,"001110000","100001001",1,'1'); -- (2, 0, 1, 1, 1, 2, 0, 0, 2)
sync_reset;
check_mem(3578,"001110010","100001001",1,'1'); -- (2, 0, 1, 1, 1, 2, 0, 1, 2)
sync_reset;
check_mem(3579,"001110000","100001010",6,'1'); -- (2, 0, 1, 1, 1, 2, 0, 2, 0)
sync_reset;
check_mem(3580,"001110001","100001010",6,'1'); -- (2, 0, 1, 1, 1, 2, 0, 2, 1)
sync_reset;
check_mem(3581,"001110000","100001100",1,'1'); -- (2, 0, 1, 1, 1, 2, 2, 0, 0)
sync_reset;
check_mem(3582,"001110001","100001100",1,'1'); -- (2, 0, 1, 1, 1, 2, 2, 0, 1)
sync_reset;
check_mem(3583,"001110010","100001100",1,'1'); -- (2, 0, 1, 1, 1, 2, 2, 1, 0)
sync_reset;
check_mem(3584,"001110010","100001101",1,'1'); -- (2, 0, 1, 1, 1, 2, 2, 1, 2)
sync_reset;
check_mem(3585,"001110001","100001110",1,'1'); -- (2, 0, 1, 1, 1, 2, 2, 2, 1)
sync_reset;
check_mem(3586,"001100000","100010000",8,'1'); -- (2, 0, 1, 1, 2, 0, 0, 0, 0)
sync_reset;
check_mem(3587,"001100001","100010000",5,'1'); -- (2, 0, 1, 1, 2, 0, 0, 0, 1)
sync_reset;
check_mem(3588,"001100010","100010000",8,'1'); -- (2, 0, 1, 1, 2, 0, 0, 1, 0)
sync_reset;
check_mem(3589,"001100001","100010010",5,'1'); -- (2, 0, 1, 1, 2, 0, 0, 2, 1)
sync_reset;
check_mem(3590,"001100100","100010000",1,'1'); -- (2, 0, 1, 1, 2, 0, 1, 0, 0)
sync_reset;
check_mem(3591,"001100100","100010010",1,'1'); -- (2, 0, 1, 1, 2, 0, 1, 2, 0)
sync_reset;
check_mem(3592,"001100101","100010010",1,'1'); -- (2, 0, 1, 1, 2, 0, 1, 2, 1)
sync_reset;
check_mem(3593,"001100001","100010100",5,'1'); -- (2, 0, 1, 1, 2, 0, 2, 0, 1)
sync_reset;
check_mem(3594,"001100010","100010100",8,'1'); -- (2, 0, 1, 1, 2, 0, 2, 1, 0)
sync_reset;
check_mem(3595,"001100011","100010100",5,'1'); -- (2, 0, 1, 1, 2, 0, 2, 1, 1)
sync_reset;
check_mem(3596,"001101000","100010000",8,'1'); -- (2, 0, 1, 1, 2, 1, 0, 0, 0)
sync_reset;
check_mem(3597,"001101000","100010010",8,'1'); -- (2, 0, 1, 1, 2, 1, 0, 2, 0)
sync_reset;
check_mem(3598,"001101100","100010010",1,'1'); -- (2, 0, 1, 1, 2, 1, 1, 2, 0)
sync_reset;
check_mem(3599,"001101000","100010100",8,'1'); -- (2, 0, 1, 1, 2, 1, 2, 0, 0)
sync_reset;
check_mem(3600,"001101010","100010100",8,'1'); -- (2, 0, 1, 1, 2, 1, 2, 1, 0)
sync_reset;
check_mem(3601,"001100001","100011000",1,'1'); -- (2, 0, 1, 1, 2, 2, 0, 0, 1)
sync_reset;
check_mem(3602,"001100010","100011000",8,'1'); -- (2, 0, 1, 1, 2, 2, 0, 1, 0)
sync_reset;
check_mem(3603,"001100011","100011000",6,'1'); -- (2, 0, 1, 1, 2, 2, 0, 1, 1)
sync_reset;
check_mem(3604,"001100100","100011000",8,'1'); -- (2, 0, 1, 1, 2, 2, 1, 0, 0)
sync_reset;
check_mem(3605,"001100101","100011000",7,'1'); -- (2, 0, 1, 1, 2, 2, 1, 0, 1)
sync_reset;
check_mem(3606,"001100110","100011000",8,'1'); -- (2, 0, 1, 1, 2, 2, 1, 1, 0)
sync_reset;
check_mem(3607,"001100101","100011010",1,'1'); -- (2, 0, 1, 1, 2, 2, 1, 2, 1)
sync_reset;
check_mem(3608,"001100011","100011100",1,'1'); -- (2, 0, 1, 1, 2, 2, 2, 1, 1)
sync_reset;
check_mem(3609,"001000001","100100000",5,'1'); -- (2, 0, 1, 2, 0, 0, 0, 0, 1)
sync_reset;
check_mem(3610,"001000010","100100000",6,'1'); -- (2, 0, 1, 2, 0, 0, 0, 1, 0)
sync_reset;
check_mem(3611,"001000011","100100000",6,'1'); -- (2, 0, 1, 2, 0, 0, 0, 1, 1)
sync_reset;
check_mem(3612,"001000100","100100000",4,'1'); -- (2, 0, 1, 2, 0, 0, 1, 0, 0)
sync_reset;
check_mem(3613,"001000101","100100000",1,'1'); -- (2, 0, 1, 2, 0, 0, 1, 0, 1)
sync_reset;
check_mem(3614,"001000110","100100000",1,'1'); -- (2, 0, 1, 2, 0, 0, 1, 1, 0)
sync_reset;
check_mem(3615,"001000110","100100001",4,'1'); -- (2, 0, 1, 2, 0, 0, 1, 1, 2)
sync_reset;
check_mem(3616,"001000101","100100010",1,'1'); -- (2, 0, 1, 2, 0, 0, 1, 2, 1)
sync_reset;
check_mem(3617,"001001000","100100000",6,'1'); -- (2, 0, 1, 2, 0, 1, 0, 0, 0)
sync_reset;
check_mem(3618,"001001010","100100000",6,'1'); -- (2, 0, 1, 2, 0, 1, 0, 1, 0)
sync_reset;
check_mem(3619,"001001010","100100001",1,'1'); -- (2, 0, 1, 2, 0, 1, 0, 1, 2)
sync_reset;
check_mem(3620,"001001100","100100000",1,'1'); -- (2, 0, 1, 2, 0, 1, 1, 0, 0)
sync_reset;
check_mem(3621,"001001100","100100001",4,'1'); -- (2, 0, 1, 2, 0, 1, 1, 0, 2)
sync_reset;
check_mem(3622,"001001110","100100001",4,'1'); -- (2, 0, 1, 2, 0, 1, 1, 1, 2)
sync_reset;
check_mem(3623,"001001100","100100010",1,'1'); -- (2, 0, 1, 2, 0, 1, 1, 2, 0)
sync_reset;
check_mem(3624,"001000011","100101000",6,'1'); -- (2, 0, 1, 2, 0, 2, 0, 1, 1)
sync_reset;
check_mem(3625,"001000101","100101000",4,'1'); -- (2, 0, 1, 2, 0, 2, 1, 0, 1)
sync_reset;
check_mem(3626,"001000110","100101000",4,'1'); -- (2, 0, 1, 2, 0, 2, 1, 1, 0)
sync_reset;
check_mem(3627,"001010000","100100000",6,'1'); -- (2, 0, 1, 2, 1, 0, 0, 0, 0)
sync_reset;
check_mem(3628,"001010001","100100000",6,'1'); -- (2, 0, 1, 2, 1, 0, 0, 0, 1)
sync_reset;
check_mem(3629,"001010010","100100000",6,'1'); -- (2, 0, 1, 2, 1, 0, 0, 1, 0)
sync_reset;
check_mem(3630,"001010010","100100001",1,'1'); -- (2, 0, 1, 2, 1, 0, 0, 1, 2)
sync_reset;
check_mem(3631,"001010001","100100010",5,'1'); -- (2, 0, 1, 2, 1, 0, 0, 2, 1)
sync_reset;
check_mem(3632,"001011000","100100000",6,'1'); -- (2, 0, 1, 2, 1, 1, 0, 0, 0)
sync_reset;
check_mem(3633,"001011000","100100001",6,'1'); -- (2, 0, 1, 2, 1, 1, 0, 0, 2)
sync_reset;
check_mem(3634,"001011010","100100001",6,'1'); -- (2, 0, 1, 2, 1, 1, 0, 1, 2)
sync_reset;
check_mem(3635,"001011000","100100010",6,'1'); -- (2, 0, 1, 2, 1, 1, 0, 2, 0)
sync_reset;
check_mem(3636,"001010001","100101000",6,'1'); -- (2, 0, 1, 2, 1, 2, 0, 0, 1)
sync_reset;
check_mem(3637,"001010010","100101000",1,'1'); -- (2, 0, 1, 2, 1, 2, 0, 1, 0)
sync_reset;
check_mem(3638,"001010011","100101000",6,'1'); -- (2, 0, 1, 2, 1, 2, 0, 1, 1)
sync_reset;
check_mem(3639,"001000011","100110000",5,'1'); -- (2, 0, 1, 2, 2, 0, 0, 1, 1)
sync_reset;
check_mem(3640,"001000101","100110000",5,'1'); -- (2, 0, 1, 2, 2, 0, 1, 0, 1)
sync_reset;
check_mem(3641,"001000110","100110000",8,'1'); -- (2, 0, 1, 2, 2, 0, 1, 1, 0)
sync_reset;
check_mem(3642,"001001010","100110000",8,'1'); -- (2, 0, 1, 2, 2, 1, 0, 1, 0)
sync_reset;
check_mem(3643,"001001100","100110000",8,'1'); -- (2, 0, 1, 2, 2, 1, 1, 0, 0)
sync_reset;
check_mem(3644,"001001110","100110000",8,'1'); -- (2, 0, 1, 2, 2, 1, 1, 1, 0)
sync_reset;
check_mem(3645,"000000011","101000000",1,'1'); -- (2, 0, 2, 0, 0, 0, 0, 1, 1)
sync_reset;
check_mem(3646,"000000101","101000000",7,'1'); -- (2, 0, 2, 0, 0, 0, 1, 0, 1)
sync_reset;
check_mem(3647,"000000110","101000000",1,'1'); -- (2, 0, 2, 0, 0, 0, 1, 1, 0)
sync_reset;
check_mem(3648,"000001001","101000000",1,'1'); -- (2, 0, 2, 0, 0, 1, 0, 0, 1)
sync_reset;
check_mem(3649,"000001010","101000000",1,'1'); -- (2, 0, 2, 0, 0, 1, 0, 1, 0)
sync_reset;
check_mem(3650,"000001011","101000000",1,'1'); -- (2, 0, 2, 0, 0, 1, 0, 1, 1)
sync_reset;
check_mem(3651,"000001100","101000000",1,'1'); -- (2, 0, 2, 0, 0, 1, 1, 0, 0)
sync_reset;
check_mem(3652,"000001101","101000000",1,'1'); -- (2, 0, 2, 0, 0, 1, 1, 0, 1)
sync_reset;
check_mem(3653,"000001110","101000000",1,'1'); -- (2, 0, 2, 0, 0, 1, 1, 1, 0)
sync_reset;
check_mem(3654,"000001110","101000001",1,'1'); -- (2, 0, 2, 0, 0, 1, 1, 1, 2)
sync_reset;
check_mem(3655,"000001101","101000010",1,'1'); -- (2, 0, 2, 0, 0, 1, 1, 2, 1)
sync_reset;
check_mem(3656,"000001011","101000100",1,'1'); -- (2, 0, 2, 0, 0, 1, 2, 1, 1)
sync_reset;
check_mem(3657,"000010001","101000000",1,'1'); -- (2, 0, 2, 0, 1, 0, 0, 0, 1)
sync_reset;
check_mem(3658,"000010010","101000000",1,'1'); -- (2, 0, 2, 0, 1, 0, 0, 1, 0)
sync_reset;
check_mem(3659,"000010011","101000000",1,'1'); -- (2, 0, 2, 0, 1, 0, 0, 1, 1)
sync_reset;
check_mem(3660,"000010100","101000000",1,'1'); -- (2, 0, 2, 0, 1, 0, 1, 0, 0)
sync_reset;
check_mem(3661,"000010101","101000000",1,'1'); -- (2, 0, 2, 0, 1, 0, 1, 0, 1)
sync_reset;
check_mem(3662,"000010110","101000000",1,'1'); -- (2, 0, 2, 0, 1, 0, 1, 1, 0)
sync_reset;
check_mem(3663,"000010110","101000001",1,'1'); -- (2, 0, 2, 0, 1, 0, 1, 1, 2)
sync_reset;
check_mem(3664,"000010101","101000010",1,'1'); -- (2, 0, 2, 0, 1, 0, 1, 2, 1)
sync_reset;
check_mem(3665,"000010011","101000100",1,'1'); -- (2, 0, 2, 0, 1, 0, 2, 1, 1)
sync_reset;
check_mem(3666,"000011000","101000000",1,'1'); -- (2, 0, 2, 0, 1, 1, 0, 0, 0)
sync_reset;
check_mem(3667,"000011001","101000000",1,'1'); -- (2, 0, 2, 0, 1, 1, 0, 0, 1)
sync_reset;
check_mem(3668,"000011010","101000000",1,'1'); -- (2, 0, 2, 0, 1, 1, 0, 1, 0)
sync_reset;
check_mem(3669,"000011010","101000001",1,'1'); -- (2, 0, 2, 0, 1, 1, 0, 1, 2)
sync_reset;
check_mem(3670,"000011001","101000010",3,'1'); -- (2, 0, 2, 0, 1, 1, 0, 2, 1)
sync_reset;
check_mem(3671,"000011100","101000000",1,'1'); -- (2, 0, 2, 0, 1, 1, 1, 0, 0)
sync_reset;
check_mem(3672,"000011100","101000001",1,'1'); -- (2, 0, 2, 0, 1, 1, 1, 0, 2)
sync_reset;
check_mem(3673,"000011110","101000001",1,'1'); -- (2, 0, 2, 0, 1, 1, 1, 1, 2)
sync_reset;
check_mem(3674,"000011100","101000010",3,'1'); -- (2, 0, 2, 0, 1, 1, 1, 2, 0)
sync_reset;
check_mem(3675,"000011101","101000010",1,'1'); -- (2, 0, 2, 0, 1, 1, 1, 2, 1)
sync_reset;
check_mem(3676,"000011001","101000100",3,'1'); -- (2, 0, 2, 0, 1, 1, 2, 0, 1)
sync_reset;
check_mem(3677,"000011010","101000100",1,'1'); -- (2, 0, 2, 0, 1, 1, 2, 1, 0)
sync_reset;
check_mem(3678,"000011011","101000100",1,'1'); -- (2, 0, 2, 0, 1, 1, 2, 1, 1)
sync_reset;
check_mem(3679,"000010011","101001000",1,'1'); -- (2, 0, 2, 0, 1, 2, 0, 1, 1)
sync_reset;
check_mem(3680,"000010101","101001000",7,'1'); -- (2, 0, 2, 0, 1, 2, 1, 0, 1)
sync_reset;
check_mem(3681,"000010110","101001000",1,'1'); -- (2, 0, 2, 0, 1, 2, 1, 1, 0)
sync_reset;
check_mem(3682,"000001011","101010000",6,'1'); -- (2, 0, 2, 0, 2, 1, 0, 1, 1)
sync_reset;
check_mem(3683,"000001101","101010000",7,'1'); -- (2, 0, 2, 0, 2, 1, 1, 0, 1)
sync_reset;
check_mem(3684,"000001110","101010000",8,'1'); -- (2, 0, 2, 0, 2, 1, 1, 1, 0)
sync_reset;
check_mem(3685,"000100001","101000000",1,'1'); -- (2, 0, 2, 1, 0, 0, 0, 0, 1)
sync_reset;
check_mem(3686,"000100010","101000000",1,'1'); -- (2, 0, 2, 1, 0, 0, 0, 1, 0)
sync_reset;
check_mem(3687,"000100011","101000000",1,'1'); -- (2, 0, 2, 1, 0, 0, 0, 1, 1)
sync_reset;
check_mem(3688,"000100100","101000000",1,'1'); -- (2, 0, 2, 1, 0, 0, 1, 0, 0)
sync_reset;
check_mem(3689,"000100101","101000000",1,'1'); -- (2, 0, 2, 1, 0, 0, 1, 0, 1)
sync_reset;
check_mem(3690,"000100110","101000000",1,'1'); -- (2, 0, 2, 1, 0, 0, 1, 1, 0)
sync_reset;
check_mem(3691,"000100110","101000001",1,'1'); -- (2, 0, 2, 1, 0, 0, 1, 1, 2)
sync_reset;
check_mem(3692,"000100101","101000010",1,'1'); -- (2, 0, 2, 1, 0, 0, 1, 2, 1)
sync_reset;
check_mem(3693,"000100011","101000100",1,'1'); -- (2, 0, 2, 1, 0, 0, 2, 1, 1)
sync_reset;
check_mem(3694,"000101000","101000000",4,'1'); -- (2, 0, 2, 1, 0, 1, 0, 0, 0)
sync_reset;
check_mem(3695,"000101001","101000000",1,'1'); -- (2, 0, 2, 1, 0, 1, 0, 0, 1)
sync_reset;
check_mem(3696,"000101010","101000000",1,'1'); -- (2, 0, 2, 1, 0, 1, 0, 1, 0)
sync_reset;
check_mem(3697,"000101010","101000001",4,'1'); -- (2, 0, 2, 1, 0, 1, 0, 1, 2)
sync_reset;
check_mem(3698,"000101001","101000010",4,'1'); -- (2, 0, 2, 1, 0, 1, 0, 2, 1)
sync_reset;
check_mem(3699,"000101100","101000000",1,'1'); -- (2, 0, 2, 1, 0, 1, 1, 0, 0)
sync_reset;
check_mem(3700,"000101100","101000001",4,'1'); -- (2, 0, 2, 1, 0, 1, 1, 0, 2)
sync_reset;
check_mem(3701,"000101110","101000001",1,'1'); -- (2, 0, 2, 1, 0, 1, 1, 1, 2)
sync_reset;
check_mem(3702,"000101100","101000010",4,'1'); -- (2, 0, 2, 1, 0, 1, 1, 2, 0)
sync_reset;
check_mem(3703,"000101101","101000010",1,'1'); -- (2, 0, 2, 1, 0, 1, 1, 2, 1)
sync_reset;
check_mem(3704,"000101001","101000100",4,'1'); -- (2, 0, 2, 1, 0, 1, 2, 0, 1)
sync_reset;
check_mem(3705,"000101010","101000100",4,'1'); -- (2, 0, 2, 1, 0, 1, 2, 1, 0)
sync_reset;
check_mem(3706,"000101011","101000100",1,'1'); -- (2, 0, 2, 1, 0, 1, 2, 1, 1)
sync_reset;
check_mem(3707,"000100011","101001000",1,'1'); -- (2, 0, 2, 1, 0, 2, 0, 1, 1)
sync_reset;
check_mem(3708,"000100101","101001000",7,'1'); -- (2, 0, 2, 1, 0, 2, 1, 0, 1)
sync_reset;
check_mem(3709,"000100110","101001000",8,'1'); -- (2, 0, 2, 1, 0, 2, 1, 1, 0)
sync_reset;
check_mem(3710,"000110000","101000000",1,'1'); -- (2, 0, 2, 1, 1, 0, 0, 0, 0)
sync_reset;
check_mem(3711,"000110001","101000000",1,'1'); -- (2, 0, 2, 1, 1, 0, 0, 0, 1)
sync_reset;
check_mem(3712,"000110010","101000000",1,'1'); -- (2, 0, 2, 1, 1, 0, 0, 1, 0)
sync_reset;
check_mem(3713,"000110010","101000001",1,'1'); -- (2, 0, 2, 1, 1, 0, 0, 1, 2)
sync_reset;
check_mem(3714,"000110001","101000010",5,'1'); -- (2, 0, 2, 1, 1, 0, 0, 2, 1)
sync_reset;
check_mem(3715,"000110100","101000000",1,'1'); -- (2, 0, 2, 1, 1, 0, 1, 0, 0)
sync_reset;
check_mem(3716,"000110100","101000001",5,'1'); -- (2, 0, 2, 1, 1, 0, 1, 0, 2)
sync_reset;
check_mem(3717,"000110110","101000001",1,'1'); -- (2, 0, 2, 1, 1, 0, 1, 1, 2)
sync_reset;
check_mem(3718,"000110100","101000010",5,'1'); -- (2, 0, 2, 1, 1, 0, 1, 2, 0)
sync_reset;
check_mem(3719,"000110101","101000010",1,'1'); -- (2, 0, 2, 1, 1, 0, 1, 2, 1)
sync_reset;
check_mem(3720,"000110001","101000100",1,'1'); -- (2, 0, 2, 1, 1, 0, 2, 0, 1)
sync_reset;
check_mem(3721,"000110010","101000100",1,'1'); -- (2, 0, 2, 1, 1, 0, 2, 1, 0)
sync_reset;
check_mem(3722,"000110011","101000100",1,'1'); -- (2, 0, 2, 1, 1, 0, 2, 1, 1)
sync_reset;
check_mem(3723,"000110001","101001000",1,'1'); -- (2, 0, 2, 1, 1, 2, 0, 0, 1)
sync_reset;
check_mem(3724,"000110010","101001000",1,'1'); -- (2, 0, 2, 1, 1, 2, 0, 1, 0)
sync_reset;
check_mem(3725,"000110011","101001000",1,'1'); -- (2, 0, 2, 1, 1, 2, 0, 1, 1)
sync_reset;
check_mem(3726,"000110100","101001000",1,'1'); -- (2, 0, 2, 1, 1, 2, 1, 0, 0)
sync_reset;
check_mem(3727,"000110101","101001000",1,'1'); -- (2, 0, 2, 1, 1, 2, 1, 0, 1)
sync_reset;
check_mem(3728,"000110110","101001000",1,'1'); -- (2, 0, 2, 1, 1, 2, 1, 1, 0)
sync_reset;
check_mem(3729,"000110101","101001010",1,'1'); -- (2, 0, 2, 1, 1, 2, 1, 2, 1)
sync_reset;
check_mem(3730,"000110011","101001100",1,'1'); -- (2, 0, 2, 1, 1, 2, 2, 1, 1)
sync_reset;
check_mem(3731,"000100011","101010000",6,'1'); -- (2, 0, 2, 1, 2, 0, 0, 1, 1)
sync_reset;
check_mem(3732,"000100101","101010000",7,'1'); -- (2, 0, 2, 1, 2, 0, 1, 0, 1)
sync_reset;
check_mem(3733,"000100110","101010000",8,'1'); -- (2, 0, 2, 1, 2, 0, 1, 1, 0)
sync_reset;
check_mem(3734,"000101001","101010000",1,'1'); -- (2, 0, 2, 1, 2, 1, 0, 0, 1)
sync_reset;
check_mem(3735,"000101010","101010000",1,'1'); -- (2, 0, 2, 1, 2, 1, 0, 1, 0)
sync_reset;
check_mem(3736,"000101011","101010000",1,'1'); -- (2, 0, 2, 1, 2, 1, 0, 1, 1)
sync_reset;
check_mem(3737,"000101100","101010000",1,'1'); -- (2, 0, 2, 1, 2, 1, 1, 0, 0)
sync_reset;
check_mem(3738,"000101101","101010000",1,'1'); -- (2, 0, 2, 1, 2, 1, 1, 0, 1)
sync_reset;
check_mem(3739,"000101110","101010000",1,'1'); -- (2, 0, 2, 1, 2, 1, 1, 1, 0)
sync_reset;
check_mem(3740,"000101101","101010010",1,'1'); -- (2, 0, 2, 1, 2, 1, 1, 2, 1)
sync_reset;
check_mem(3741,"000001011","101100000",6,'1'); -- (2, 0, 2, 2, 0, 1, 0, 1, 1)
sync_reset;
check_mem(3742,"000001101","101100000",7,'1'); -- (2, 0, 2, 2, 0, 1, 1, 0, 1)
sync_reset;
check_mem(3743,"000001110","101100000",1,'1'); -- (2, 0, 2, 2, 0, 1, 1, 1, 0)
sync_reset;
check_mem(3744,"000010011","101100000",1,'1'); -- (2, 0, 2, 2, 1, 0, 0, 1, 1)
sync_reset;
check_mem(3745,"000010101","101100000",7,'1'); -- (2, 0, 2, 2, 1, 0, 1, 0, 1)
sync_reset;
check_mem(3746,"000010110","101100000",1,'1'); -- (2, 0, 2, 2, 1, 0, 1, 1, 0)
sync_reset;
check_mem(3747,"000011001","101100000",1,'1'); -- (2, 0, 2, 2, 1, 1, 0, 0, 1)
sync_reset;
check_mem(3748,"000011010","101100000",1,'1'); -- (2, 0, 2, 2, 1, 1, 0, 1, 0)
sync_reset;
check_mem(3749,"000011011","101100000",1,'1'); -- (2, 0, 2, 2, 1, 1, 0, 1, 1)
sync_reset;
check_mem(3750,"000011100","101100000",1,'1'); -- (2, 0, 2, 2, 1, 1, 1, 0, 0)
sync_reset;
check_mem(3751,"000011101","101100000",1,'1'); -- (2, 0, 2, 2, 1, 1, 1, 0, 1)
sync_reset;
check_mem(3752,"000011110","101100000",1,'1'); -- (2, 0, 2, 2, 1, 1, 1, 1, 0)
sync_reset;
check_mem(3753,"000011110","101100001",1,'1'); -- (2, 0, 2, 2, 1, 1, 1, 1, 2)
sync_reset;
check_mem(3754,"000011101","101100010",1,'1'); -- (2, 0, 2, 2, 1, 1, 1, 2, 1)
sync_reset;
check_mem(3755,"010000000","100000000",3,'1'); -- (2, 1, 0, 0, 0, 0, 0, 0, 0)
sync_reset;
check_mem(3756,"010000001","100000000",4,'1'); -- (2, 1, 0, 0, 0, 0, 0, 0, 1)
sync_reset;
check_mem(3757,"010000010","100000000",4,'1'); -- (2, 1, 0, 0, 0, 0, 0, 1, 0)
sync_reset;
check_mem(3758,"010000010","100000001",4,'1'); -- (2, 1, 0, 0, 0, 0, 0, 1, 2)
sync_reset;
check_mem(3759,"010000001","100000010",2,'1'); -- (2, 1, 0, 0, 0, 0, 0, 2, 1)
sync_reset;
check_mem(3760,"010000100","100000000",4,'1'); -- (2, 1, 0, 0, 0, 0, 1, 0, 0)
sync_reset;
check_mem(3761,"010000100","100000001",4,'1'); -- (2, 1, 0, 0, 0, 0, 1, 0, 2)
sync_reset;
check_mem(3762,"010000110","100000001",4,'1'); -- (2, 1, 0, 0, 0, 0, 1, 1, 2)
sync_reset;
check_mem(3763,"010000100","100000010",2,'1'); -- (2, 1, 0, 0, 0, 0, 1, 2, 0)
sync_reset;
check_mem(3764,"010000101","100000010",2,'1'); -- (2, 1, 0, 0, 0, 0, 1, 2, 1)
sync_reset;
check_mem(3765,"010000001","100000100",3,'1'); -- (2, 1, 0, 0, 0, 0, 2, 0, 1)
sync_reset;
check_mem(3766,"010000010","100000100",4,'1'); -- (2, 1, 0, 0, 0, 0, 2, 1, 0)
sync_reset;
check_mem(3767,"010000011","100000100",3,'1'); -- (2, 1, 0, 0, 0, 0, 2, 1, 1)
sync_reset;
check_mem(3768,"010001000","100000000",6,'1'); -- (2, 1, 0, 0, 0, 1, 0, 0, 0)
sync_reset;
check_mem(3769,"010001000","100000001",4,'1'); -- (2, 1, 0, 0, 0, 1, 0, 0, 2)
sync_reset;
check_mem(3770,"010001010","100000001",4,'1'); -- (2, 1, 0, 0, 0, 1, 0, 1, 2)
sync_reset;
check_mem(3771,"010001000","100000010",3,'1'); -- (2, 1, 0, 0, 0, 1, 0, 2, 0)
sync_reset;
check_mem(3772,"010001001","100000010",2,'1'); -- (2, 1, 0, 0, 0, 1, 0, 2, 1)
sync_reset;
check_mem(3773,"010001100","100000001",4,'1'); -- (2, 1, 0, 0, 0, 1, 1, 0, 2)
sync_reset;
check_mem(3774,"010001100","100000010",2,'1'); -- (2, 1, 0, 0, 0, 1, 1, 2, 0)
sync_reset;
check_mem(3775,"010001100","100000011",4,'1'); -- (2, 1, 0, 0, 0, 1, 1, 2, 2)
sync_reset;
check_mem(3776,"010001000","100000100",2,'1'); -- (2, 1, 0, 0, 0, 1, 2, 0, 0)
sync_reset;
check_mem(3777,"010001001","100000100",2,'1'); -- (2, 1, 0, 0, 0, 1, 2, 0, 1)
sync_reset;
check_mem(3778,"010001010","100000100",3,'1'); -- (2, 1, 0, 0, 0, 1, 2, 1, 0)
sync_reset;
check_mem(3779,"010001010","100000101",4,'1'); -- (2, 1, 0, 0, 0, 1, 2, 1, 2)
sync_reset;
check_mem(3780,"010001001","100000110",2,'1'); -- (2, 1, 0, 0, 0, 1, 2, 2, 1)
sync_reset;
check_mem(3781,"010000001","100001000",7,'1'); -- (2, 1, 0, 0, 0, 2, 0, 0, 1)
sync_reset;
check_mem(3782,"010000010","100001000",4,'1'); -- (2, 1, 0, 0, 0, 2, 0, 1, 0)
sync_reset;
check_mem(3783,"010000011","100001000",2,'1'); -- (2, 1, 0, 0, 0, 2, 0, 1, 1)
sync_reset;
check_mem(3784,"010000100","100001000",4,'1'); -- (2, 1, 0, 0, 0, 2, 1, 0, 0)
sync_reset;
check_mem(3785,"010000101","100001000",7,'1'); -- (2, 1, 0, 0, 0, 2, 1, 0, 1)
sync_reset;
check_mem(3786,"010000110","100001000",2,'1'); -- (2, 1, 0, 0, 0, 2, 1, 1, 0)
sync_reset;
check_mem(3787,"010000110","100001001",4,'1'); -- (2, 1, 0, 0, 0, 2, 1, 1, 2)
sync_reset;
check_mem(3788,"010000101","100001010",2,'1'); -- (2, 1, 0, 0, 0, 2, 1, 2, 1)
sync_reset;
check_mem(3789,"010000011","100001100",4,'1'); -- (2, 1, 0, 0, 0, 2, 2, 1, 1)
sync_reset;
check_mem(3790,"010010000","100000000",7,'1'); -- (2, 1, 0, 0, 1, 0, 0, 0, 0)
sync_reset;
check_mem(3791,"010010000","100000001",2,'1'); -- (2, 1, 0, 0, 1, 0, 0, 0, 2)
sync_reset;
check_mem(3792,"010010000","100000010",3,'1'); -- (2, 1, 0, 0, 1, 0, 0, 2, 0)
sync_reset;
check_mem(3793,"010010001","100000010",2,'1'); -- (2, 1, 0, 0, 1, 0, 0, 2, 1)
sync_reset;
check_mem(3794,"010010100","100000001",2,'1'); -- (2, 1, 0, 0, 1, 0, 1, 0, 2)
sync_reset;
check_mem(3795,"010010100","100000010",2,'1'); -- (2, 1, 0, 0, 1, 0, 1, 2, 0)
sync_reset;
check_mem(3796,"010010100","100000011",2,'1'); -- (2, 1, 0, 0, 1, 0, 1, 2, 2)
sync_reset;
check_mem(3797,"010010000","100000100",3,'1'); -- (2, 1, 0, 0, 1, 0, 2, 0, 0)
sync_reset;
check_mem(3798,"010010001","100000100",3,'1'); -- (2, 1, 0, 0, 1, 0, 2, 0, 1)
sync_reset;
check_mem(3799,"010010001","100000110",3,'1'); -- (2, 1, 0, 0, 1, 0, 2, 2, 1)
sync_reset;
check_mem(3800,"010011000","100000001",2,'1'); -- (2, 1, 0, 0, 1, 1, 0, 0, 2)
sync_reset;
check_mem(3801,"010011000","100000010",3,'1'); -- (2, 1, 0, 0, 1, 1, 0, 2, 0)
sync_reset;
check_mem(3802,"010011000","100000011",3,'1'); -- (2, 1, 0, 0, 1, 1, 0, 2, 2)
sync_reset;
check_mem(3803,"010011100","100000011",2,'1'); -- (2, 1, 0, 0, 1, 1, 1, 2, 2)
sync_reset;
check_mem(3804,"010011000","100000100",3,'1'); -- (2, 1, 0, 0, 1, 1, 2, 0, 0)
sync_reset;
check_mem(3805,"010011000","100000101",3,'1'); -- (2, 1, 0, 0, 1, 1, 2, 0, 2)
sync_reset;
check_mem(3806,"010011000","100000110",3,'1'); -- (2, 1, 0, 0, 1, 1, 2, 2, 0)
sync_reset;
check_mem(3807,"010011001","100000110",3,'1'); -- (2, 1, 0, 0, 1, 1, 2, 2, 1)
sync_reset;
check_mem(3808,"010010000","100001000",2,'1'); -- (2, 1, 0, 0, 1, 2, 0, 0, 0)
sync_reset;
check_mem(3809,"010010001","100001000",7,'1'); -- (2, 1, 0, 0, 1, 2, 0, 0, 1)
sync_reset;
check_mem(3810,"010010001","100001010",2,'1'); -- (2, 1, 0, 0, 1, 2, 0, 2, 1)
sync_reset;
check_mem(3811,"010010100","100001000",2,'1'); -- (2, 1, 0, 0, 1, 2, 1, 0, 0)
sync_reset;
check_mem(3812,"010010100","100001001",2,'1'); -- (2, 1, 0, 0, 1, 2, 1, 0, 2)
sync_reset;
check_mem(3813,"010010100","100001010",2,'1'); -- (2, 1, 0, 0, 1, 2, 1, 2, 0)
sync_reset;
check_mem(3814,"010010101","100001010",2,'1'); -- (2, 1, 0, 0, 1, 2, 1, 2, 1)
sync_reset;
check_mem(3815,"010010001","100001100",7,'1'); -- (2, 1, 0, 0, 1, 2, 2, 0, 1)
sync_reset;
check_mem(3816,"010000001","100010000",2,'1'); -- (2, 1, 0, 0, 2, 0, 0, 0, 1)
sync_reset;
check_mem(3817,"010000010","100010000",2,'1'); -- (2, 1, 0, 0, 2, 0, 0, 1, 0)
sync_reset;
check_mem(3818,"010000011","100010000",6,'1'); -- (2, 1, 0, 0, 2, 0, 0, 1, 1)
sync_reset;
check_mem(3819,"010000100","100010000",8,'1'); -- (2, 1, 0, 0, 2, 0, 1, 0, 0)
sync_reset;
check_mem(3820,"010000101","100010000",7,'1'); -- (2, 1, 0, 0, 2, 0, 1, 0, 1)
sync_reset;
check_mem(3821,"010000110","100010000",8,'1'); -- (2, 1, 0, 0, 2, 0, 1, 1, 0)
sync_reset;
check_mem(3822,"010000101","100010010",2,'1'); -- (2, 1, 0, 0, 2, 0, 1, 2, 1)
sync_reset;
check_mem(3823,"010000011","100010100",2,'1'); -- (2, 1, 0, 0, 2, 0, 2, 1, 1)
sync_reset;
check_mem(3824,"010001000","100010000",8,'1'); -- (2, 1, 0, 0, 2, 1, 0, 0, 0)
sync_reset;
check_mem(3825,"010001001","100010000",2,'1'); -- (2, 1, 0, 0, 2, 1, 0, 0, 1)
sync_reset;
check_mem(3826,"010001010","100010000",2,'1'); -- (2, 1, 0, 0, 2, 1, 0, 1, 0)
sync_reset;
check_mem(3827,"010001001","100010010",2,'1'); -- (2, 1, 0, 0, 2, 1, 0, 2, 1)
sync_reset;
check_mem(3828,"010001100","100010000",8,'1'); -- (2, 1, 0, 0, 2, 1, 1, 0, 0)
sync_reset;
check_mem(3829,"010001100","100010010",8,'1'); -- (2, 1, 0, 0, 2, 1, 1, 2, 0)
sync_reset;
check_mem(3830,"010001101","100010010",2,'1'); -- (2, 1, 0, 0, 2, 1, 1, 2, 1)
sync_reset;
check_mem(3831,"010001001","100010100",2,'1'); -- (2, 1, 0, 0, 2, 1, 2, 0, 1)
sync_reset;
check_mem(3832,"010001010","100010100",2,'1'); -- (2, 1, 0, 0, 2, 1, 2, 1, 0)
sync_reset;
check_mem(3833,"010001011","100010100",2,'1'); -- (2, 1, 0, 0, 2, 1, 2, 1, 1)
sync_reset;
check_mem(3834,"010000011","100011000",6,'1'); -- (2, 1, 0, 0, 2, 2, 0, 1, 1)
sync_reset;
check_mem(3835,"010000101","100011000",7,'1'); -- (2, 1, 0, 0, 2, 2, 1, 0, 1)
sync_reset;
check_mem(3836,"010000110","100011000",8,'1'); -- (2, 1, 0, 0, 2, 2, 1, 1, 0)
sync_reset;
check_mem(3837,"010100000","100000000",4,'1'); -- (2, 1, 0, 1, 0, 0, 0, 0, 0)
sync_reset;
check_mem(3838,"010100000","100000001",4,'1'); -- (2, 1, 0, 1, 0, 0, 0, 0, 2)
sync_reset;
check_mem(3839,"010100010","100000001",4,'1'); -- (2, 1, 0, 1, 0, 0, 0, 1, 2)
sync_reset;
check_mem(3840,"010100000","100000010",4,'1'); -- (2, 1, 0, 1, 0, 0, 0, 2, 0)
sync_reset;
check_mem(3841,"010100001","100000010",2,'1'); -- (2, 1, 0, 1, 0, 0, 0, 2, 1)
sync_reset;
check_mem(3842,"010100100","100000001",2,'1'); -- (2, 1, 0, 1, 0, 0, 1, 0, 2)
sync_reset;
check_mem(3843,"010100100","100000010",2,'1'); -- (2, 1, 0, 1, 0, 0, 1, 2, 0)
sync_reset;
check_mem(3844,"010100100","100000011",4,'1'); -- (2, 1, 0, 1, 0, 0, 1, 2, 2)
sync_reset;
check_mem(3845,"010100000","100000100",4,'1'); -- (2, 1, 0, 1, 0, 0, 2, 0, 0)
sync_reset;
check_mem(3846,"010100001","100000100",4,'1'); -- (2, 1, 0, 1, 0, 0, 2, 0, 1)
sync_reset;
check_mem(3847,"010100010","100000100",4,'1'); -- (2, 1, 0, 1, 0, 0, 2, 1, 0)
sync_reset;
check_mem(3848,"010100010","100000101",4,'1'); -- (2, 1, 0, 1, 0, 0, 2, 1, 2)
sync_reset;
check_mem(3849,"010100001","100000110",5,'1'); -- (2, 1, 0, 1, 0, 0, 2, 2, 1)
sync_reset;
check_mem(3850,"010101000","100000001",4,'1'); -- (2, 1, 0, 1, 0, 1, 0, 0, 2)
sync_reset;
check_mem(3851,"010101000","100000010",4,'1'); -- (2, 1, 0, 1, 0, 1, 0, 2, 0)
sync_reset;
check_mem(3852,"010101000","100000011",4,'1'); -- (2, 1, 0, 1, 0, 1, 0, 2, 2)
sync_reset;
check_mem(3853,"010101100","100000011",4,'1'); -- (2, 1, 0, 1, 0, 1, 1, 2, 2)
sync_reset;
check_mem(3854,"010101000","100000100",4,'1'); -- (2, 1, 0, 1, 0, 1, 2, 0, 0)
sync_reset;
check_mem(3855,"010101000","100000101",4,'1'); -- (2, 1, 0, 1, 0, 1, 2, 0, 2)
sync_reset;
check_mem(3856,"010101010","100000101",4,'1'); -- (2, 1, 0, 1, 0, 1, 2, 1, 2)
sync_reset;
check_mem(3857,"010101000","100000110",4,'1'); -- (2, 1, 0, 1, 0, 1, 2, 2, 0)
sync_reset;
check_mem(3858,"010101001","100000110",2,'1'); -- (2, 1, 0, 1, 0, 1, 2, 2, 1)
sync_reset;
check_mem(3859,"010100000","100001000",2,'1'); -- (2, 1, 0, 1, 0, 2, 0, 0, 0)
sync_reset;
check_mem(3860,"010100001","100001000",4,'1'); -- (2, 1, 0, 1, 0, 2, 0, 0, 1)
sync_reset;
check_mem(3861,"010100010","100001000",4,'1'); -- (2, 1, 0, 1, 0, 2, 0, 1, 0)
sync_reset;
check_mem(3862,"010100010","100001001",4,'1'); -- (2, 1, 0, 1, 0, 2, 0, 1, 2)
sync_reset;
check_mem(3863,"010100001","100001010",2,'1'); -- (2, 1, 0, 1, 0, 2, 0, 2, 1)
sync_reset;
check_mem(3864,"010100100","100001000",8,'1'); -- (2, 1, 0, 1, 0, 2, 1, 0, 0)
sync_reset;
check_mem(3865,"010100100","100001001",2,'1'); -- (2, 1, 0, 1, 0, 2, 1, 0, 2)
sync_reset;
check_mem(3866,"010100110","100001001",2,'1'); -- (2, 1, 0, 1, 0, 2, 1, 1, 2)
sync_reset;
check_mem(3867,"010100100","100001010",2,'1'); -- (2, 1, 0, 1, 0, 2, 1, 2, 0)
sync_reset;
check_mem(3868,"010100101","100001010",2,'1'); -- (2, 1, 0, 1, 0, 2, 1, 2, 1)
sync_reset;
check_mem(3869,"010100001","100001100",2,'1'); -- (2, 1, 0, 1, 0, 2, 2, 0, 1)
sync_reset;
check_mem(3870,"010100010","100001100",4,'1'); -- (2, 1, 0, 1, 0, 2, 2, 1, 0)
sync_reset;
check_mem(3871,"010100011","100001100",4,'1'); -- (2, 1, 0, 1, 0, 2, 2, 1, 1)
sync_reset;
check_mem(3872,"010110000","100000001",2,'1'); -- (2, 1, 0, 1, 1, 0, 0, 0, 2)
sync_reset;
check_mem(3873,"010110000","100000010",5,'1'); -- (2, 1, 0, 1, 1, 0, 0, 2, 0)
sync_reset;
check_mem(3874,"010110000","100000011",5,'1'); -- (2, 1, 0, 1, 1, 0, 0, 2, 2)
sync_reset;
check_mem(3875,"010110100","100000011",2,'1'); -- (2, 1, 0, 1, 1, 0, 1, 2, 2)
sync_reset;
check_mem(3876,"010110000","100000100",2,'1'); -- (2, 1, 0, 1, 1, 0, 2, 0, 0)
sync_reset;
check_mem(3877,"010110000","100000101",5,'1'); -- (2, 1, 0, 1, 1, 0, 2, 0, 2)
sync_reset;
check_mem(3878,"010110000","100000110",5,'1'); -- (2, 1, 0, 1, 1, 0, 2, 2, 0)
sync_reset;
check_mem(3879,"010110001","100000110",5,'1'); -- (2, 1, 0, 1, 1, 0, 2, 2, 1)
sync_reset;
check_mem(3880,"010110000","100001000",7,'1'); -- (2, 1, 0, 1, 1, 2, 0, 0, 0)
sync_reset;
check_mem(3881,"010110000","100001001",2,'1'); -- (2, 1, 0, 1, 1, 2, 0, 0, 2)
sync_reset;
check_mem(3882,"010110000","100001010",2,'1'); -- (2, 1, 0, 1, 1, 2, 0, 2, 0)
sync_reset;
check_mem(3883,"010110001","100001010",2,'1'); -- (2, 1, 0, 1, 1, 2, 0, 2, 1)
sync_reset;
check_mem(3884,"010110100","100001001",2,'1'); -- (2, 1, 0, 1, 1, 2, 1, 0, 2)
sync_reset;
check_mem(3885,"010110100","100001010",2,'1'); -- (2, 1, 0, 1, 1, 2, 1, 2, 0)
sync_reset;
check_mem(3886,"010110100","100001011",2,'1'); -- (2, 1, 0, 1, 1, 2, 1, 2, 2)
sync_reset;
check_mem(3887,"010110000","100001100",7,'1'); -- (2, 1, 0, 1, 1, 2, 2, 0, 0)
sync_reset;
check_mem(3888,"010110001","100001100",7,'1'); -- (2, 1, 0, 1, 1, 2, 2, 0, 1)
sync_reset;
check_mem(3889,"010110001","100001110",2,'1'); -- (2, 1, 0, 1, 1, 2, 2, 2, 1)
sync_reset;
check_mem(3890,"010100000","100010000",8,'1'); -- (2, 1, 0, 1, 2, 0, 0, 0, 0)
sync_reset;
check_mem(3891,"010100001","100010000",2,'1'); -- (2, 1, 0, 1, 2, 0, 0, 0, 1)
sync_reset;
check_mem(3892,"010100010","100010000",2,'1'); -- (2, 1, 0, 1, 2, 0, 0, 1, 0)
sync_reset;
check_mem(3893,"010100001","100010010",2,'1'); -- (2, 1, 0, 1, 2, 0, 0, 2, 1)
sync_reset;
check_mem(3894,"010100100","100010000",8,'1'); -- (2, 1, 0, 1, 2, 0, 1, 0, 0)
sync_reset;
check_mem(3895,"010100100","100010010",8,'1'); -- (2, 1, 0, 1, 2, 0, 1, 2, 0)
sync_reset;
check_mem(3896,"010100101","100010010",2,'1'); -- (2, 1, 0, 1, 2, 0, 1, 2, 1)
sync_reset;
check_mem(3897,"010100001","100010100",2,'1'); -- (2, 1, 0, 1, 2, 0, 2, 0, 1)
sync_reset;
check_mem(3898,"010100010","100010100",2,'1'); -- (2, 1, 0, 1, 2, 0, 2, 1, 0)
sync_reset;
check_mem(3899,"010100011","100010100",2,'1'); -- (2, 1, 0, 1, 2, 0, 2, 1, 1)
sync_reset;
check_mem(3900,"010101000","100010000",2,'1'); -- (2, 1, 0, 1, 2, 1, 0, 0, 0)
sync_reset;
check_mem(3901,"010101000","100010010",8,'1'); -- (2, 1, 0, 1, 2, 1, 0, 2, 0)
sync_reset;
check_mem(3902,"010101001","100010010",2,'1'); -- (2, 1, 0, 1, 2, 1, 0, 2, 1)
sync_reset;
check_mem(3903,"010101100","100010010",8,'1'); -- (2, 1, 0, 1, 2, 1, 1, 2, 0)
sync_reset;
check_mem(3904,"010101000","100010100",2,'1'); -- (2, 1, 0, 1, 2, 1, 2, 0, 0)
sync_reset;
check_mem(3905,"010101001","100010100",2,'1'); -- (2, 1, 0, 1, 2, 1, 2, 0, 1)
sync_reset;
check_mem(3906,"010101010","100010100",2,'1'); -- (2, 1, 0, 1, 2, 1, 2, 1, 0)
sync_reset;
check_mem(3907,"010101001","100010110",2,'1'); -- (2, 1, 0, 1, 2, 1, 2, 2, 1)
sync_reset;
check_mem(3908,"010100001","100011000",2,'1'); -- (2, 1, 0, 1, 2, 2, 0, 0, 1)
sync_reset;
check_mem(3909,"010100010","100011000",8,'1'); -- (2, 1, 0, 1, 2, 2, 0, 1, 0)
sync_reset;
check_mem(3910,"010100011","100011000",6,'1'); -- (2, 1, 0, 1, 2, 2, 0, 1, 1)
sync_reset;
check_mem(3911,"010100100","100011000",8,'1'); -- (2, 1, 0, 1, 2, 2, 1, 0, 0)
sync_reset;
check_mem(3912,"010100101","100011000",7,'1'); -- (2, 1, 0, 1, 2, 2, 1, 0, 1)
sync_reset;
check_mem(3913,"010100110","100011000",8,'1'); -- (2, 1, 0, 1, 2, 2, 1, 1, 0)
sync_reset;
check_mem(3914,"010100101","100011010",2,'1'); -- (2, 1, 0, 1, 2, 2, 1, 2, 1)
sync_reset;
check_mem(3915,"010100011","100011100",2,'1'); -- (2, 1, 0, 1, 2, 2, 2, 1, 1)
sync_reset;
check_mem(3916,"010000001","100100000",6,'1'); -- (2, 1, 0, 2, 0, 0, 0, 0, 1)
sync_reset;
check_mem(3917,"010000010","100100000",4,'1'); -- (2, 1, 0, 2, 0, 0, 0, 1, 0)
sync_reset;
check_mem(3918,"010000011","100100000",6,'1'); -- (2, 1, 0, 2, 0, 0, 0, 1, 1)
sync_reset;
check_mem(3919,"010000100","100100000",4,'1'); -- (2, 1, 0, 2, 0, 0, 1, 0, 0)
sync_reset;
check_mem(3920,"010000101","100100000",2,'1'); -- (2, 1, 0, 2, 0, 0, 1, 0, 1)
sync_reset;
check_mem(3921,"010000110","100100000",2,'1'); -- (2, 1, 0, 2, 0, 0, 1, 1, 0)
sync_reset;
check_mem(3922,"010000110","100100001",4,'1'); -- (2, 1, 0, 2, 0, 0, 1, 1, 2)
sync_reset;
check_mem(3923,"010000101","100100010",2,'1'); -- (2, 1, 0, 2, 0, 0, 1, 2, 1)
sync_reset;
check_mem(3924,"010001000","100100000",6,'1'); -- (2, 1, 0, 2, 0, 1, 0, 0, 0)
sync_reset;
check_mem(3925,"010001001","100100000",6,'1'); -- (2, 1, 0, 2, 0, 1, 0, 0, 1)
sync_reset;
check_mem(3926,"010001010","100100000",4,'1'); -- (2, 1, 0, 2, 0, 1, 0, 1, 0)
sync_reset;
check_mem(3927,"010001010","100100001",4,'1'); -- (2, 1, 0, 2, 0, 1, 0, 1, 2)
sync_reset;
check_mem(3928,"010001001","100100010",2,'1'); -- (2, 1, 0, 2, 0, 1, 0, 2, 1)
sync_reset;
check_mem(3929,"010001100","100100000",2,'1'); -- (2, 1, 0, 2, 0, 1, 1, 0, 0)
sync_reset;
check_mem(3930,"010001100","100100001",4,'1'); -- (2, 1, 0, 2, 0, 1, 1, 0, 2)
sync_reset;
check_mem(3931,"010001110","100100001",4,'1'); -- (2, 1, 0, 2, 0, 1, 1, 1, 2)
sync_reset;
check_mem(3932,"010001100","100100010",2,'1'); -- (2, 1, 0, 2, 0, 1, 1, 2, 0)
sync_reset;
check_mem(3933,"010001101","100100010",2,'1'); -- (2, 1, 0, 2, 0, 1, 1, 2, 1)
sync_reset;
check_mem(3934,"010000011","100101000",4,'1'); -- (2, 1, 0, 2, 0, 2, 0, 1, 1)
sync_reset;
check_mem(3935,"010000101","100101000",4,'1'); -- (2, 1, 0, 2, 0, 2, 1, 0, 1)
sync_reset;
check_mem(3936,"010000110","100101000",4,'1'); -- (2, 1, 0, 2, 0, 2, 1, 1, 0)
sync_reset;
check_mem(3937,"010010000","100100000",6,'1'); -- (2, 1, 0, 2, 1, 0, 0, 0, 0)
sync_reset;
check_mem(3938,"010010001","100100000",6,'1'); -- (2, 1, 0, 2, 1, 0, 0, 0, 1)
sync_reset;
check_mem(3939,"010010001","100100010",6,'1'); -- (2, 1, 0, 2, 1, 0, 0, 2, 1)
sync_reset;
check_mem(3940,"010010100","100100000",2,'1'); -- (2, 1, 0, 2, 1, 0, 1, 0, 0)
sync_reset;
check_mem(3941,"010010100","100100001",2,'1'); -- (2, 1, 0, 2, 1, 0, 1, 0, 2)
sync_reset;
check_mem(3942,"010010100","100100010",2,'1'); -- (2, 1, 0, 2, 1, 0, 1, 2, 0)
sync_reset;
check_mem(3943,"010010101","100100010",2,'1'); -- (2, 1, 0, 2, 1, 0, 1, 2, 1)
sync_reset;
check_mem(3944,"010011000","100100000",6,'1'); -- (2, 1, 0, 2, 1, 1, 0, 0, 0)
sync_reset;
check_mem(3945,"010011000","100100001",6,'1'); -- (2, 1, 0, 2, 1, 1, 0, 0, 2)
sync_reset;
check_mem(3946,"010011000","100100010",6,'1'); -- (2, 1, 0, 2, 1, 1, 0, 2, 0)
sync_reset;
check_mem(3947,"010011001","100100010",6,'1'); -- (2, 1, 0, 2, 1, 1, 0, 2, 1)
sync_reset;
check_mem(3948,"010011100","100100001",2,'1'); -- (2, 1, 0, 2, 1, 1, 1, 0, 2)
sync_reset;
check_mem(3949,"010011100","100100010",2,'1'); -- (2, 1, 0, 2, 1, 1, 1, 2, 0)
sync_reset;
check_mem(3950,"010011100","100100011",2,'1'); -- (2, 1, 0, 2, 1, 1, 1, 2, 2)
sync_reset;
check_mem(3951,"010010001","100101000",6,'1'); -- (2, 1, 0, 2, 1, 2, 0, 0, 1)
sync_reset;
check_mem(3952,"010010100","100101000",2,'1'); -- (2, 1, 0, 2, 1, 2, 1, 0, 0)
sync_reset;
check_mem(3953,"010010101","100101000",2,'1'); -- (2, 1, 0, 2, 1, 2, 1, 0, 1)
sync_reset;
check_mem(3954,"010010101","100101010",2,'1'); -- (2, 1, 0, 2, 1, 2, 1, 2, 1)
sync_reset;
check_mem(3955,"010000011","100110000",6,'1'); -- (2, 1, 0, 2, 2, 0, 0, 1, 1)
sync_reset;
check_mem(3956,"010000101","100110000",5,'1'); -- (2, 1, 0, 2, 2, 0, 1, 0, 1)
sync_reset;
check_mem(3957,"010000110","100110000",8,'1'); -- (2, 1, 0, 2, 2, 0, 1, 1, 0)
sync_reset;
check_mem(3958,"010001001","100110000",2,'1'); -- (2, 1, 0, 2, 2, 1, 0, 0, 1)
sync_reset;
check_mem(3959,"010001010","100110000",2,'1'); -- (2, 1, 0, 2, 2, 1, 0, 1, 0)
sync_reset;
check_mem(3960,"010001011","100110000",6,'1'); -- (2, 1, 0, 2, 2, 1, 0, 1, 1)
sync_reset;
check_mem(3961,"010001100","100110000",8,'1'); -- (2, 1, 0, 2, 2, 1, 1, 0, 0)
sync_reset;
check_mem(3962,"010001101","100110000",2,'1'); -- (2, 1, 0, 2, 2, 1, 1, 0, 1)
sync_reset;
check_mem(3963,"010001110","100110000",8,'1'); -- (2, 1, 0, 2, 2, 1, 1, 1, 0)
sync_reset;
check_mem(3964,"010001101","100110010",2,'1'); -- (2, 1, 0, 2, 2, 1, 1, 2, 1)
sync_reset;
check_mem(3965,"011000000","100000000",3,'1'); -- (2, 1, 1, 0, 0, 0, 0, 0, 0)
sync_reset;
check_mem(3966,"011000000","100000001",4,'1'); -- (2, 1, 1, 0, 0, 0, 0, 0, 2)
sync_reset;
check_mem(3967,"011000010","100000001",4,'1'); -- (2, 1, 1, 0, 0, 0, 0, 1, 2)
sync_reset;
check_mem(3968,"011000000","100000010",6,'1'); -- (2, 1, 1, 0, 0, 0, 0, 2, 0)
sync_reset;
check_mem(3969,"011000001","100000010",5,'1'); -- (2, 1, 1, 0, 0, 0, 0, 2, 1)
sync_reset;
check_mem(3970,"011000100","100000001",4,'1'); -- (2, 1, 1, 0, 0, 0, 1, 0, 2)
sync_reset;
check_mem(3971,"011000100","100000010",4,'1'); -- (2, 1, 1, 0, 0, 0, 1, 2, 0)
sync_reset;
check_mem(3972,"011000100","100000011",4,'1'); -- (2, 1, 1, 0, 0, 0, 1, 2, 2)
sync_reset;
check_mem(3973,"011000000","100000100",3,'1'); -- (2, 1, 1, 0, 0, 0, 2, 0, 0)
sync_reset;
check_mem(3974,"011000001","100000100",3,'1'); -- (2, 1, 1, 0, 0, 0, 2, 0, 1)
sync_reset;
check_mem(3975,"011000010","100000100",3,'1'); -- (2, 1, 1, 0, 0, 0, 2, 1, 0)
sync_reset;
check_mem(3976,"011000010","100000101",4,'1'); -- (2, 1, 1, 0, 0, 0, 2, 1, 2)
sync_reset;
check_mem(3977,"011000001","100000110",5,'1'); -- (2, 1, 1, 0, 0, 0, 2, 2, 1)
sync_reset;
check_mem(3978,"011001000","100000001",3,'1'); -- (2, 1, 1, 0, 0, 1, 0, 0, 2)
sync_reset;
check_mem(3979,"011001000","100000010",8,'1'); -- (2, 1, 1, 0, 0, 1, 0, 2, 0)
sync_reset;
check_mem(3980,"011001000","100000011",3,'1'); -- (2, 1, 1, 0, 0, 1, 0, 2, 2)
sync_reset;
check_mem(3981,"011001100","100000011",4,'1'); -- (2, 1, 1, 0, 0, 1, 1, 2, 2)
sync_reset;
check_mem(3982,"011001000","100000100",3,'1'); -- (2, 1, 1, 0, 0, 1, 2, 0, 0)
sync_reset;
check_mem(3983,"011001000","100000101",3,'1'); -- (2, 1, 1, 0, 0, 1, 2, 0, 2)
sync_reset;
check_mem(3984,"011001010","100000101",3,'1'); -- (2, 1, 1, 0, 0, 1, 2, 1, 2)
sync_reset;
check_mem(3985,"011001000","100000110",8,'1'); -- (2, 1, 1, 0, 0, 1, 2, 2, 0)
sync_reset;
check_mem(3986,"011000000","100001000",4,'1'); -- (2, 1, 1, 0, 0, 2, 0, 0, 0)
sync_reset;
check_mem(3987,"011000001","100001000",3,'1'); -- (2, 1, 1, 0, 0, 2, 0, 0, 1)
sync_reset;
check_mem(3988,"011000010","100001000",4,'1'); -- (2, 1, 1, 0, 0, 2, 0, 1, 0)
sync_reset;
check_mem(3989,"011000010","100001001",4,'1'); -- (2, 1, 1, 0, 0, 2, 0, 1, 2)
sync_reset;
check_mem(3990,"011000001","100001010",3,'1'); -- (2, 1, 1, 0, 0, 2, 0, 2, 1)
sync_reset;
check_mem(3991,"011000100","100001000",4,'1'); -- (2, 1, 1, 0, 0, 2, 1, 0, 0)
sync_reset;
check_mem(3992,"011000100","100001001",4,'1'); -- (2, 1, 1, 0, 0, 2, 1, 0, 2)
sync_reset;
check_mem(3993,"011000110","100001001",4,'1'); -- (2, 1, 1, 0, 0, 2, 1, 1, 2)
sync_reset;
check_mem(3994,"011000100","100001010",4,'1'); -- (2, 1, 1, 0, 0, 2, 1, 2, 0)
sync_reset;
check_mem(3995,"011000101","100001010",4,'1'); -- (2, 1, 1, 0, 0, 2, 1, 2, 1)
sync_reset;
check_mem(3996,"011000001","100001100",3,'1'); -- (2, 1, 1, 0, 0, 2, 2, 0, 1)
sync_reset;
check_mem(3997,"011000010","100001100",4,'1'); -- (2, 1, 1, 0, 0, 2, 2, 1, 0)
sync_reset;
check_mem(3998,"011000011","100001100",3,'1'); -- (2, 1, 1, 0, 0, 2, 2, 1, 1)
sync_reset;
check_mem(3999,"011010000","100000001",3,'1'); -- (2, 1, 1, 0, 1, 0, 0, 0, 2)
sync_reset;
check_mem(4000,"011010000","100000010",6,'1'); -- (2, 1, 1, 0, 1, 0, 0, 2, 0)
sync_reset;
check_mem(4001,"011010000","100000011",6,'1'); -- (2, 1, 1, 0, 1, 0, 0, 2, 2)
sync_reset;
check_mem(4002,"011010000","100000100",3,'1'); -- (2, 1, 1, 0, 1, 0, 2, 0, 0)
sync_reset;
check_mem(4003,"011010000","100000101",7,'1'); -- (2, 1, 1, 0, 1, 0, 2, 0, 2)
sync_reset;
check_mem(4004,"011010000","100000110",3,'1'); -- (2, 1, 1, 0, 1, 0, 2, 2, 0)
sync_reset;
check_mem(4005,"011010001","100000110",3,'1'); -- (2, 1, 1, 0, 1, 0, 2, 2, 1)
sync_reset;
check_mem(4006,"011011000","100000011",6,'1'); -- (2, 1, 1, 0, 1, 1, 0, 2, 2)
sync_reset;
check_mem(4007,"011011000","100000101",3,'1'); -- (2, 1, 1, 0, 1, 1, 2, 0, 2)
sync_reset;
check_mem(4008,"011011000","100000110",3,'1'); -- (2, 1, 1, 0, 1, 1, 2, 2, 0)
sync_reset;
check_mem(4009,"011010000","100001000",3,'1'); -- (2, 1, 1, 0, 1, 2, 0, 0, 0)
sync_reset;
check_mem(4010,"011010000","100001001",3,'1'); -- (2, 1, 1, 0, 1, 2, 0, 0, 2)
sync_reset;
check_mem(4011,"011010000","100001010",6,'1'); -- (2, 1, 1, 0, 1, 2, 0, 2, 0)
sync_reset;
check_mem(4012,"011010001","100001010",6,'1'); -- (2, 1, 1, 0, 1, 2, 0, 2, 1)
sync_reset;
check_mem(4013,"011010000","100001100",7,'1'); -- (2, 1, 1, 0, 1, 2, 2, 0, 0)
sync_reset;
check_mem(4014,"011010001","100001100",3,'1'); -- (2, 1, 1, 0, 1, 2, 2, 0, 1)
sync_reset;
check_mem(4015,"011010001","100001110",3,'1'); -- (2, 1, 1, 0, 1, 2, 2, 2, 1)
sync_reset;
check_mem(4016,"011000000","100010000",8,'1'); -- (2, 1, 1, 0, 2, 0, 0, 0, 0)
sync_reset;
check_mem(4017,"011000001","100010000",5,'1'); -- (2, 1, 1, 0, 2, 0, 0, 0, 1)
sync_reset;
check_mem(4018,"011000010","100010000",3,'1'); -- (2, 1, 1, 0, 2, 0, 0, 1, 0)
sync_reset;
check_mem(4019,"011000001","100010010",5,'1'); -- (2, 1, 1, 0, 2, 0, 0, 2, 1)
sync_reset;
check_mem(4020,"011000100","100010000",3,'1'); -- (2, 1, 1, 0, 2, 0, 1, 0, 0)
sync_reset;
check_mem(4021,"011000100","100010010",8,'1'); -- (2, 1, 1, 0, 2, 0, 1, 2, 0)
sync_reset;
check_mem(4022,"011000101","100010010",5,'1'); -- (2, 1, 1, 0, 2, 0, 1, 2, 1)
sync_reset;
check_mem(4023,"011000001","100010100",5,'1'); -- (2, 1, 1, 0, 2, 0, 2, 0, 1)
sync_reset;
check_mem(4024,"011000010","100010100",3,'1'); -- (2, 1, 1, 0, 2, 0, 2, 1, 0)
sync_reset;
check_mem(4025,"011000011","100010100",3,'1'); -- (2, 1, 1, 0, 2, 0, 2, 1, 1)
sync_reset;
check_mem(4026,"011001000","100010000",8,'1'); -- (2, 1, 1, 0, 2, 1, 0, 0, 0)
sync_reset;
check_mem(4027,"011001000","100010010",8,'1'); -- (2, 1, 1, 0, 2, 1, 0, 2, 0)
sync_reset;
check_mem(4028,"011001100","100010010",8,'1'); -- (2, 1, 1, 0, 2, 1, 1, 2, 0)
sync_reset;
check_mem(4029,"011001000","100010100",8,'1'); -- (2, 1, 1, 0, 2, 1, 2, 0, 0)
sync_reset;
check_mem(4030,"011001010","100010100",3,'1'); -- (2, 1, 1, 0, 2, 1, 2, 1, 0)
sync_reset;
check_mem(4031,"011000001","100011000",3,'1'); -- (2, 1, 1, 0, 2, 2, 0, 0, 1)
sync_reset;
check_mem(4032,"011000010","100011000",3,'1'); -- (2, 1, 1, 0, 2, 2, 0, 1, 0)
sync_reset;
check_mem(4033,"011000011","100011000",3,'1'); -- (2, 1, 1, 0, 2, 2, 0, 1, 1)
sync_reset;
check_mem(4034,"011000100","100011000",3,'1'); -- (2, 1, 1, 0, 2, 2, 1, 0, 0)
sync_reset;
check_mem(4035,"011000101","100011000",3,'1'); -- (2, 1, 1, 0, 2, 2, 1, 0, 1)
sync_reset;
check_mem(4036,"011000110","100011000",3,'1'); -- (2, 1, 1, 0, 2, 2, 1, 1, 0)
sync_reset;
check_mem(4037,"011000101","100011010",3,'1'); -- (2, 1, 1, 0, 2, 2, 1, 2, 1)
sync_reset;
check_mem(4038,"011000011","100011100",3,'1'); -- (2, 1, 1, 0, 2, 2, 2, 1, 1)
sync_reset;
check_mem(4039,"011100000","100000001",4,'1'); -- (2, 1, 1, 1, 0, 0, 0, 0, 2)
sync_reset;
check_mem(4040,"011100000","100000010",8,'1'); -- (2, 1, 1, 1, 0, 0, 0, 2, 0)
sync_reset;
check_mem(4041,"011100000","100000011",4,'1'); -- (2, 1, 1, 1, 0, 0, 0, 2, 2)
sync_reset;
check_mem(4042,"011100100","100000011",4,'1'); -- (2, 1, 1, 1, 0, 0, 1, 2, 2)
sync_reset;
check_mem(4043,"011100000","100000100",8,'1'); -- (2, 1, 1, 1, 0, 0, 2, 0, 0)
sync_reset;
check_mem(4044,"011100000","100000101",4,'1'); -- (2, 1, 1, 1, 0, 0, 2, 0, 2)
sync_reset;
check_mem(4045,"011100010","100000101",4,'1'); -- (2, 1, 1, 1, 0, 0, 2, 1, 2)
sync_reset;
check_mem(4046,"011100000","100000110",8,'1'); -- (2, 1, 1, 1, 0, 0, 2, 2, 0)
sync_reset;
check_mem(4047,"011100001","100000110",5,'1'); -- (2, 1, 1, 1, 0, 0, 2, 2, 1)
sync_reset;
check_mem(4048,"011101000","100000011",4,'1'); -- (2, 1, 1, 1, 0, 1, 0, 2, 2)
sync_reset;
check_mem(4049,"011101000","100000101",4,'1'); -- (2, 1, 1, 1, 0, 1, 2, 0, 2)
sync_reset;
check_mem(4050,"011101000","100000110",8,'1'); -- (2, 1, 1, 1, 0, 1, 2, 2, 0)
sync_reset;
check_mem(4051,"011100000","100001000",4,'1'); -- (2, 1, 1, 1, 0, 2, 0, 0, 0)
sync_reset;
check_mem(4052,"011100000","100001001",4,'1'); -- (2, 1, 1, 1, 0, 2, 0, 0, 2)
sync_reset;
check_mem(4053,"011100010","100001001",4,'1'); -- (2, 1, 1, 1, 0, 2, 0, 1, 2)
sync_reset;
check_mem(4054,"011100000","100001010",4,'1'); -- (2, 1, 1, 1, 0, 2, 0, 2, 0)
sync_reset;
check_mem(4055,"011100001","100001010",4,'1'); -- (2, 1, 1, 1, 0, 2, 0, 2, 1)
sync_reset;
check_mem(4056,"011100100","100001001",4,'1'); -- (2, 1, 1, 1, 0, 2, 1, 0, 2)
sync_reset;
check_mem(4057,"011100100","100001010",4,'1'); -- (2, 1, 1, 1, 0, 2, 1, 2, 0)
sync_reset;
check_mem(4058,"011100100","100001011",4,'1'); -- (2, 1, 1, 1, 0, 2, 1, 2, 2)
sync_reset;
check_mem(4059,"011100000","100001100",4,'1'); -- (2, 1, 1, 1, 0, 2, 2, 0, 0)
sync_reset;
check_mem(4060,"011100001","100001100",4,'1'); -- (2, 1, 1, 1, 0, 2, 2, 0, 1)
sync_reset;
check_mem(4061,"011100010","100001100",4,'1'); -- (2, 1, 1, 1, 0, 2, 2, 1, 0)
sync_reset;
check_mem(4062,"011100010","100001101",4,'1'); -- (2, 1, 1, 1, 0, 2, 2, 1, 2)
sync_reset;
check_mem(4063,"011100001","100001110",4,'1'); -- (2, 1, 1, 1, 0, 2, 2, 2, 1)
sync_reset;
check_mem(4064,"011110000","100000011",6,'1'); -- (2, 1, 1, 1, 1, 0, 0, 2, 2)
sync_reset;
check_mem(4065,"011110000","100000101",7,'1'); -- (2, 1, 1, 1, 1, 0, 2, 0, 2)
sync_reset;
check_mem(4066,"011110000","100000110",8,'1'); -- (2, 1, 1, 1, 1, 0, 2, 2, 0)
sync_reset;
check_mem(4067,"011110000","100001001",6,'1'); -- (2, 1, 1, 1, 1, 2, 0, 0, 2)
sync_reset;
check_mem(4068,"011110000","100001010",6,'1'); -- (2, 1, 1, 1, 1, 2, 0, 2, 0)
sync_reset;
check_mem(4069,"011110000","100001011",6,'1'); -- (2, 1, 1, 1, 1, 2, 0, 2, 2)
sync_reset;
check_mem(4070,"011110000","100001100",7,'1'); -- (2, 1, 1, 1, 1, 2, 2, 0, 0)
sync_reset;
check_mem(4071,"011110000","100001101",7,'1'); -- (2, 1, 1, 1, 1, 2, 2, 0, 2)
sync_reset;
check_mem(4072,"011110000","100001110",8,'1'); -- (2, 1, 1, 1, 1, 2, 2, 2, 0)
sync_reset;
check_mem(4073,"011100000","100010000",8,'1'); -- (2, 1, 1, 1, 2, 0, 0, 0, 0)
sync_reset;
check_mem(4074,"011100000","100010010",8,'1'); -- (2, 1, 1, 1, 2, 0, 0, 2, 0)
sync_reset;
check_mem(4075,"011100001","100010010",5,'1'); -- (2, 1, 1, 1, 2, 0, 0, 2, 1)
sync_reset;
check_mem(4076,"011100100","100010010",8,'1'); -- (2, 1, 1, 1, 2, 0, 1, 2, 0)
sync_reset;
check_mem(4077,"011100000","100010100",8,'1'); -- (2, 1, 1, 1, 2, 0, 2, 0, 0)
sync_reset;
check_mem(4078,"011100001","100010100",5,'1'); -- (2, 1, 1, 1, 2, 0, 2, 0, 1)
sync_reset;
check_mem(4079,"011100010","100010100",8,'1'); -- (2, 1, 1, 1, 2, 0, 2, 1, 0)
sync_reset;
check_mem(4080,"011100001","100010110",5,'1'); -- (2, 1, 1, 1, 2, 0, 2, 2, 1)
sync_reset;
check_mem(4081,"011101000","100010010",8,'1'); -- (2, 1, 1, 1, 2, 1, 0, 2, 0)
sync_reset;
check_mem(4082,"011101000","100010100",8,'1'); -- (2, 1, 1, 1, 2, 1, 2, 0, 0)
sync_reset;
check_mem(4083,"011101000","100010110",8,'1'); -- (2, 1, 1, 1, 2, 1, 2, 2, 0)
sync_reset;
check_mem(4084,"011100000","100011000",8,'1'); -- (2, 1, 1, 1, 2, 2, 0, 0, 0)
sync_reset;
check_mem(4085,"011100001","100011000",6,'1'); -- (2, 1, 1, 1, 2, 2, 0, 0, 1)
sync_reset;
check_mem(4086,"011100010","100011000",8,'1'); -- (2, 1, 1, 1, 2, 2, 0, 1, 0)
sync_reset;
check_mem(4087,"011100001","100011010",6,'1'); -- (2, 1, 1, 1, 2, 2, 0, 2, 1)
sync_reset;
check_mem(4088,"011100100","100011000",8,'1'); -- (2, 1, 1, 1, 2, 2, 1, 0, 0)
sync_reset;
check_mem(4089,"011100100","100011010",8,'1'); -- (2, 1, 1, 1, 2, 2, 1, 2, 0)
sync_reset;
check_mem(4090,"011100001","100011100",7,'1'); -- (2, 1, 1, 1, 2, 2, 2, 0, 1)
sync_reset;
check_mem(4091,"011100010","100011100",8,'1'); -- (2, 1, 1, 1, 2, 2, 2, 1, 0)
sync_reset;
check_mem(4092,"011000000","100100000",4,'1'); -- (2, 1, 1, 2, 0, 0, 0, 0, 0)
sync_reset;
check_mem(4093,"011000001","100100000",5,'1'); -- (2, 1, 1, 2, 0, 0, 0, 0, 1)
sync_reset;
check_mem(4094,"011000010","100100000",4,'1'); -- (2, 1, 1, 2, 0, 0, 0, 1, 0)
sync_reset;
check_mem(4095,"011000010","100100001",4,'1'); -- (2, 1, 1, 2, 0, 0, 0, 1, 2)
sync_reset;
check_mem(4096,"011000001","100100010",5,'1'); -- (2, 1, 1, 2, 0, 0, 0, 2, 1)
sync_reset;
check_mem(4097,"011000100","100100000",4,'1'); -- (2, 1, 1, 2, 0, 0, 1, 0, 0)
sync_reset;
check_mem(4098,"011000100","100100001",4,'1'); -- (2, 1, 1, 2, 0, 0, 1, 0, 2)
sync_reset;
check_mem(4099,"011000110","100100001",4,'1'); -- (2, 1, 1, 2, 0, 0, 1, 1, 2)
sync_reset;
check_mem(4100,"011000100","100100010",4,'1'); -- (2, 1, 1, 2, 0, 0, 1, 2, 0)
sync_reset;
check_mem(4101,"011000101","100100010",4,'1'); -- (2, 1, 1, 2, 0, 0, 1, 2, 1)
sync_reset;
check_mem(4102,"011001000","100100000",6,'1'); -- (2, 1, 1, 2, 0, 1, 0, 0, 0)
sync_reset;
check_mem(4103,"011001000","100100001",4,'1'); -- (2, 1, 1, 2, 0, 1, 0, 0, 2)
sync_reset;
check_mem(4104,"011001010","100100001",4,'1'); -- (2, 1, 1, 2, 0, 1, 0, 1, 2)
sync_reset;
check_mem(4105,"011001000","100100010",6,'1'); -- (2, 1, 1, 2, 0, 1, 0, 2, 0)
sync_reset;
check_mem(4106,"011001100","100100001",4,'1'); -- (2, 1, 1, 2, 0, 1, 1, 0, 2)
sync_reset;
check_mem(4107,"011001100","100100010",4,'1'); -- (2, 1, 1, 2, 0, 1, 1, 2, 0)
sync_reset;
check_mem(4108,"011001100","100100011",4,'1'); -- (2, 1, 1, 2, 0, 1, 1, 2, 2)
sync_reset;
check_mem(4109,"011000001","100101000",4,'1'); -- (2, 1, 1, 2, 0, 2, 0, 0, 1)
sync_reset;
check_mem(4110,"011000010","100101000",4,'1'); -- (2, 1, 1, 2, 0, 2, 0, 1, 0)
sync_reset;
check_mem(4111,"011000011","100101000",4,'1'); -- (2, 1, 1, 2, 0, 2, 0, 1, 1)
sync_reset;
check_mem(4112,"011000100","100101000",4,'1'); -- (2, 1, 1, 2, 0, 2, 1, 0, 0)
sync_reset;
check_mem(4113,"011000101","100101000",4,'1'); -- (2, 1, 1, 2, 0, 2, 1, 0, 1)
sync_reset;
check_mem(4114,"011000110","100101000",4,'1'); -- (2, 1, 1, 2, 0, 2, 1, 1, 0)
sync_reset;
check_mem(4115,"011000110","100101001",4,'1'); -- (2, 1, 1, 2, 0, 2, 1, 1, 2)
sync_reset;
check_mem(4116,"011000101","100101010",4,'1'); -- (2, 1, 1, 2, 0, 2, 1, 2, 1)
sync_reset;
check_mem(4117,"011010000","100100000",6,'1'); -- (2, 1, 1, 2, 1, 0, 0, 0, 0)
sync_reset;
check_mem(4118,"011010000","100100001",6,'1'); -- (2, 1, 1, 2, 1, 0, 0, 0, 2)
sync_reset;
check_mem(4119,"011010000","100100010",6,'1'); -- (2, 1, 1, 2, 1, 0, 0, 2, 0)
sync_reset;
check_mem(4120,"011010001","100100010",6,'1'); -- (2, 1, 1, 2, 1, 0, 0, 2, 1)
sync_reset;
check_mem(4121,"011011000","100100001",6,'1'); -- (2, 1, 1, 2, 1, 1, 0, 0, 2)
sync_reset;
check_mem(4122,"011011000","100100010",6,'1'); -- (2, 1, 1, 2, 1, 1, 0, 2, 0)
sync_reset;
check_mem(4123,"011011000","100100011",6,'1'); -- (2, 1, 1, 2, 1, 1, 0, 2, 2)
sync_reset;
check_mem(4124,"011010000","100101000",6,'1'); -- (2, 1, 1, 2, 1, 2, 0, 0, 0)
sync_reset;
check_mem(4125,"011010001","100101000",6,'1'); -- (2, 1, 1, 2, 1, 2, 0, 0, 1)
sync_reset;
check_mem(4126,"011010001","100101010",6,'1'); -- (2, 1, 1, 2, 1, 2, 0, 2, 1)
sync_reset;
check_mem(4127,"011000001","100110000",5,'1'); -- (2, 1, 1, 2, 2, 0, 0, 0, 1)
sync_reset;
check_mem(4128,"011000010","100110000",5,'1'); -- (2, 1, 1, 2, 2, 0, 0, 1, 0)
sync_reset;
check_mem(4129,"011000011","100110000",5,'1'); -- (2, 1, 1, 2, 2, 0, 0, 1, 1)
sync_reset;
check_mem(4130,"011000100","100110000",5,'1'); -- (2, 1, 1, 2, 2, 0, 1, 0, 0)
sync_reset;
check_mem(4131,"011000101","100110000",5,'1'); -- (2, 1, 1, 2, 2, 0, 1, 0, 1)
sync_reset;
check_mem(4132,"011000110","100110000",5,'1'); -- (2, 1, 1, 2, 2, 0, 1, 1, 0)
sync_reset;
check_mem(4133,"011000101","100110010",5,'1'); -- (2, 1, 1, 2, 2, 0, 1, 2, 1)
sync_reset;
check_mem(4134,"011001000","100110000",8,'1'); -- (2, 1, 1, 2, 2, 1, 0, 0, 0)
sync_reset;
check_mem(4135,"011001010","100110000",6,'1'); -- (2, 1, 1, 2, 2, 1, 0, 1, 0)
sync_reset;
check_mem(4136,"011001100","100110000",8,'1'); -- (2, 1, 1, 2, 2, 1, 1, 0, 0)
sync_reset;
check_mem(4137,"011001100","100110010",8,'1'); -- (2, 1, 1, 2, 2, 1, 1, 2, 0)
sync_reset;
check_mem(4138,"010000001","101000000",7,'1'); -- (2, 1, 2, 0, 0, 0, 0, 0, 1)
sync_reset;
check_mem(4139,"010000010","101000000",4,'1'); -- (2, 1, 2, 0, 0, 0, 0, 1, 0)
sync_reset;
check_mem(4140,"010000011","101000000",3,'1'); -- (2, 1, 2, 0, 0, 0, 0, 1, 1)
sync_reset;
check_mem(4141,"010000100","101000000",7,'1'); -- (2, 1, 2, 0, 0, 0, 1, 0, 0)
sync_reset;
check_mem(4142,"010000101","101000000",7,'1'); -- (2, 1, 2, 0, 0, 0, 1, 0, 1)
sync_reset;
check_mem(4143,"010000110","101000000",3,'1'); -- (2, 1, 2, 0, 0, 0, 1, 1, 0)
sync_reset;
check_mem(4144,"010000110","101000001",4,'1'); -- (2, 1, 2, 0, 0, 0, 1, 1, 2)
sync_reset;
check_mem(4145,"010000101","101000010",3,'1'); -- (2, 1, 2, 0, 0, 0, 1, 2, 1)
sync_reset;
check_mem(4146,"010000011","101000100",4,'1'); -- (2, 1, 2, 0, 0, 0, 2, 1, 1)
sync_reset;
check_mem(4147,"010001000","101000000",4,'1'); -- (2, 1, 2, 0, 0, 1, 0, 0, 0)
sync_reset;
check_mem(4148,"010001001","101000000",6,'1'); -- (2, 1, 2, 0, 0, 1, 0, 0, 1)
sync_reset;
check_mem(4149,"010001010","101000000",4,'1'); -- (2, 1, 2, 0, 0, 1, 0, 1, 0)
sync_reset;
check_mem(4150,"010001010","101000001",4,'1'); -- (2, 1, 2, 0, 0, 1, 0, 1, 2)
sync_reset;
check_mem(4151,"010001001","101000010",3,'1'); -- (2, 1, 2, 0, 0, 1, 0, 2, 1)
sync_reset;
check_mem(4152,"010001100","101000000",4,'1'); -- (2, 1, 2, 0, 0, 1, 1, 0, 0)
sync_reset;
check_mem(4153,"010001100","101000001",4,'1'); -- (2, 1, 2, 0, 0, 1, 1, 0, 2)
sync_reset;
check_mem(4154,"010001110","101000001",4,'1'); -- (2, 1, 2, 0, 0, 1, 1, 1, 2)
sync_reset;
check_mem(4155,"010001100","101000010",3,'1'); -- (2, 1, 2, 0, 0, 1, 1, 2, 0)
sync_reset;
check_mem(4156,"010001101","101000010",3,'1'); -- (2, 1, 2, 0, 0, 1, 1, 2, 1)
sync_reset;
check_mem(4157,"010001001","101000100",3,'1'); -- (2, 1, 2, 0, 0, 1, 2, 0, 1)
sync_reset;
check_mem(4158,"010001010","101000100",4,'1'); -- (2, 1, 2, 0, 0, 1, 2, 1, 0)
sync_reset;
check_mem(4159,"010001011","101000100",3,'1'); -- (2, 1, 2, 0, 0, 1, 2, 1, 1)
sync_reset;
check_mem(4160,"010000011","101001000",3,'1'); -- (2, 1, 2, 0, 0, 2, 0, 1, 1)
sync_reset;
check_mem(4161,"010000101","101001000",7,'1'); -- (2, 1, 2, 0, 0, 2, 1, 0, 1)
sync_reset;
check_mem(4162,"010000110","101001000",4,'1'); -- (2, 1, 2, 0, 0, 2, 1, 1, 0)
sync_reset;
check_mem(4163,"010010000","101000000",3,'1'); -- (2, 1, 2, 0, 1, 0, 0, 0, 0)
sync_reset;
check_mem(4164,"010010001","101000000",7,'1'); -- (2, 1, 2, 0, 1, 0, 0, 0, 1)
sync_reset;
check_mem(4165,"010010001","101000010",3,'1'); -- (2, 1, 2, 0, 1, 0, 0, 2, 1)
sync_reset;
check_mem(4166,"010010100","101000000",7,'1'); -- (2, 1, 2, 0, 1, 0, 1, 0, 0)
sync_reset;
check_mem(4167,"010010100","101000001",5,'1'); -- (2, 1, 2, 0, 1, 0, 1, 0, 2)
sync_reset;
check_mem(4168,"010010100","101000010",3,'1'); -- (2, 1, 2, 0, 1, 0, 1, 2, 0)
sync_reset;
check_mem(4169,"010010101","101000010",3,'1'); -- (2, 1, 2, 0, 1, 0, 1, 2, 1)
sync_reset;
check_mem(4170,"010010001","101000100",3,'1'); -- (2, 1, 2, 0, 1, 0, 2, 0, 1)
sync_reset;
check_mem(4171,"010011000","101000000",3,'1'); -- (2, 1, 2, 0, 1, 1, 0, 0, 0)
sync_reset;
check_mem(4172,"010011000","101000001",3,'1'); -- (2, 1, 2, 0, 1, 1, 0, 0, 2)
sync_reset;
check_mem(4173,"010011000","101000010",3,'1'); -- (2, 1, 2, 0, 1, 1, 0, 2, 0)
sync_reset;
check_mem(4174,"010011001","101000010",3,'1'); -- (2, 1, 2, 0, 1, 1, 0, 2, 1)
sync_reset;
check_mem(4175,"010011100","101000001",3,'1'); -- (2, 1, 2, 0, 1, 1, 1, 0, 2)
sync_reset;
check_mem(4176,"010011100","101000010",3,'1'); -- (2, 1, 2, 0, 1, 1, 1, 2, 0)
sync_reset;
check_mem(4177,"010011100","101000011",3,'1'); -- (2, 1, 2, 0, 1, 1, 1, 2, 2)
sync_reset;
check_mem(4178,"010011000","101000100",3,'1'); -- (2, 1, 2, 0, 1, 1, 2, 0, 0)
sync_reset;
check_mem(4179,"010011001","101000100",3,'1'); -- (2, 1, 2, 0, 1, 1, 2, 0, 1)
sync_reset;
check_mem(4180,"010011001","101000110",3,'1'); -- (2, 1, 2, 0, 1, 1, 2, 2, 1)
sync_reset;
check_mem(4181,"010010001","101001000",7,'1'); -- (2, 1, 2, 0, 1, 2, 0, 0, 1)
sync_reset;
check_mem(4182,"010010100","101001000",7,'1'); -- (2, 1, 2, 0, 1, 2, 1, 0, 0)
sync_reset;
check_mem(4183,"010010101","101001000",7,'1'); -- (2, 1, 2, 0, 1, 2, 1, 0, 1)
sync_reset;
check_mem(4184,"010010101","101001010",3,'1'); -- (2, 1, 2, 0, 1, 2, 1, 2, 1)
sync_reset;
check_mem(4185,"010000011","101010000",6,'1'); -- (2, 1, 2, 0, 2, 0, 0, 1, 1)
sync_reset;
check_mem(4186,"010000101","101010000",7,'1'); -- (2, 1, 2, 0, 2, 0, 1, 0, 1)
sync_reset;
check_mem(4187,"010000110","101010000",8,'1'); -- (2, 1, 2, 0, 2, 0, 1, 1, 0)
sync_reset;
check_mem(4188,"010001001","101010000",6,'1'); -- (2, 1, 2, 0, 2, 1, 0, 0, 1)
sync_reset;
check_mem(4189,"010001010","101010000",3,'1'); -- (2, 1, 2, 0, 2, 1, 0, 1, 0)
sync_reset;
check_mem(4190,"010001011","101010000",6,'1'); -- (2, 1, 2, 0, 2, 1, 0, 1, 1)
sync_reset;
check_mem(4191,"010001100","101010000",8,'1'); -- (2, 1, 2, 0, 2, 1, 1, 0, 0)
sync_reset;
check_mem(4192,"010001101","101010000",7,'1'); -- (2, 1, 2, 0, 2, 1, 1, 0, 1)
sync_reset;
check_mem(4193,"010001110","101010000",8,'1'); -- (2, 1, 2, 0, 2, 1, 1, 1, 0)
sync_reset;
check_mem(4194,"010001101","101010010",3,'1'); -- (2, 1, 2, 0, 2, 1, 1, 2, 1)
sync_reset;
check_mem(4195,"010100000","101000000",4,'1'); -- (2, 1, 2, 1, 0, 0, 0, 0, 0)
sync_reset;
check_mem(4196,"010100001","101000000",4,'1'); -- (2, 1, 2, 1, 0, 0, 0, 0, 1)
sync_reset;
check_mem(4197,"010100010","101000000",4,'1'); -- (2, 1, 2, 1, 0, 0, 0, 1, 0)
sync_reset;
check_mem(4198,"010100010","101000001",4,'1'); -- (2, 1, 2, 1, 0, 0, 0, 1, 2)
sync_reset;
check_mem(4199,"010100001","101000010",4,'1'); -- (2, 1, 2, 1, 0, 0, 0, 2, 1)
sync_reset;
check_mem(4200,"010100100","101000000",8,'1'); -- (2, 1, 2, 1, 0, 0, 1, 0, 0)
sync_reset;
check_mem(4201,"010100100","101000001",4,'1'); -- (2, 1, 2, 1, 0, 0, 1, 0, 2)
sync_reset;
check_mem(4202,"010100110","101000001",4,'1'); -- (2, 1, 2, 1, 0, 0, 1, 1, 2)
sync_reset;
check_mem(4203,"010100100","101000010",4,'1'); -- (2, 1, 2, 1, 0, 0, 1, 2, 0)
sync_reset;
check_mem(4204,"010100101","101000010",4,'1'); -- (2, 1, 2, 1, 0, 0, 1, 2, 1)
sync_reset;
check_mem(4205,"010100001","101000100",4,'1'); -- (2, 1, 2, 1, 0, 0, 2, 0, 1)
sync_reset;
check_mem(4206,"010100010","101000100",4,'1'); -- (2, 1, 2, 1, 0, 0, 2, 1, 0)
sync_reset;
check_mem(4207,"010100011","101000100",4,'1'); -- (2, 1, 2, 1, 0, 0, 2, 1, 1)
sync_reset;
check_mem(4208,"010101000","101000000",4,'1'); -- (2, 1, 2, 1, 0, 1, 0, 0, 0)
sync_reset;
check_mem(4209,"010101000","101000001",4,'1'); -- (2, 1, 2, 1, 0, 1, 0, 0, 2)
sync_reset;
check_mem(4210,"010101010","101000001",4,'1'); -- (2, 1, 2, 1, 0, 1, 0, 1, 2)
sync_reset;
check_mem(4211,"010101000","101000010",4,'1'); -- (2, 1, 2, 1, 0, 1, 0, 2, 0)
sync_reset;
check_mem(4212,"010101001","101000010",4,'1'); -- (2, 1, 2, 1, 0, 1, 0, 2, 1)
sync_reset;
check_mem(4213,"010101100","101000001",4,'1'); -- (2, 1, 2, 1, 0, 1, 1, 0, 2)
sync_reset;
check_mem(4214,"010101100","101000010",4,'1'); -- (2, 1, 2, 1, 0, 1, 1, 2, 0)
sync_reset;
check_mem(4215,"010101100","101000011",4,'1'); -- (2, 1, 2, 1, 0, 1, 1, 2, 2)
sync_reset;
check_mem(4216,"010101000","101000100",4,'1'); -- (2, 1, 2, 1, 0, 1, 2, 0, 0)
sync_reset;
check_mem(4217,"010101001","101000100",4,'1'); -- (2, 1, 2, 1, 0, 1, 2, 0, 1)
sync_reset;
check_mem(4218,"010101010","101000100",4,'1'); -- (2, 1, 2, 1, 0, 1, 2, 1, 0)
sync_reset;
check_mem(4219,"010101010","101000101",4,'1'); -- (2, 1, 2, 1, 0, 1, 2, 1, 2)
sync_reset;
check_mem(4220,"010101001","101000110",4,'1'); -- (2, 1, 2, 1, 0, 1, 2, 2, 1)
sync_reset;
check_mem(4221,"010100001","101001000",7,'1'); -- (2, 1, 2, 1, 0, 2, 0, 0, 1)
sync_reset;
check_mem(4222,"010100010","101001000",4,'1'); -- (2, 1, 2, 1, 0, 2, 0, 1, 0)
sync_reset;
check_mem(4223,"010100011","101001000",4,'1'); -- (2, 1, 2, 1, 0, 2, 0, 1, 1)
sync_reset;
check_mem(4224,"010100100","101001000",8,'1'); -- (2, 1, 2, 1, 0, 2, 1, 0, 0)
sync_reset;
check_mem(4225,"010100101","101001000",7,'1'); -- (2, 1, 2, 1, 0, 2, 1, 0, 1)
sync_reset;
check_mem(4226,"010100110","101001000",8,'1'); -- (2, 1, 2, 1, 0, 2, 1, 1, 0)
sync_reset;
check_mem(4227,"010100101","101001010",4,'1'); -- (2, 1, 2, 1, 0, 2, 1, 2, 1)
sync_reset;
check_mem(4228,"010100011","101001100",4,'1'); -- (2, 1, 2, 1, 0, 2, 2, 1, 1)
sync_reset;
check_mem(4229,"010110000","101000000",5,'1'); -- (2, 1, 2, 1, 1, 0, 0, 0, 0)
sync_reset;
check_mem(4230,"010110000","101000001",5,'1'); -- (2, 1, 2, 1, 1, 0, 0, 0, 2)
sync_reset;
check_mem(4231,"010110000","101000010",5,'1'); -- (2, 1, 2, 1, 1, 0, 0, 2, 0)
sync_reset;
check_mem(4232,"010110001","101000010",5,'1'); -- (2, 1, 2, 1, 1, 0, 0, 2, 1)
sync_reset;
check_mem(4233,"010110100","101000001",5,'1'); -- (2, 1, 2, 1, 1, 0, 1, 0, 2)
sync_reset;
check_mem(4234,"010110100","101000010",5,'1'); -- (2, 1, 2, 1, 1, 0, 1, 2, 0)
sync_reset;
check_mem(4235,"010110100","101000011",5,'1'); -- (2, 1, 2, 1, 1, 0, 1, 2, 2)
sync_reset;
check_mem(4236,"010110000","101000100",5,'1'); -- (2, 1, 2, 1, 1, 0, 2, 0, 0)
sync_reset;
check_mem(4237,"010110001","101000100",5,'1'); -- (2, 1, 2, 1, 1, 0, 2, 0, 1)
sync_reset;
check_mem(4238,"010110001","101000110",5,'1'); -- (2, 1, 2, 1, 1, 0, 2, 2, 1)
sync_reset;
check_mem(4239,"010110000","101001000",7,'1'); -- (2, 1, 2, 1, 1, 2, 0, 0, 0)
sync_reset;
check_mem(4240,"010110001","101001000",7,'1'); -- (2, 1, 2, 1, 1, 2, 0, 0, 1)
sync_reset;
check_mem(4241,"010110001","101001010",6,'1'); -- (2, 1, 2, 1, 1, 2, 0, 2, 1)
sync_reset;
check_mem(4242,"010110100","101001000",8,'1'); -- (2, 1, 2, 1, 1, 2, 1, 0, 0)
sync_reset;
check_mem(4243,"010110100","101001010",8,'1'); -- (2, 1, 2, 1, 1, 2, 1, 2, 0)
sync_reset;
check_mem(4244,"010110001","101001100",7,'1'); -- (2, 1, 2, 1, 1, 2, 2, 0, 1)
sync_reset;
check_mem(4245,"010100001","101010000",6,'1'); -- (2, 1, 2, 1, 2, 0, 0, 0, 1)
sync_reset;
check_mem(4246,"010100010","101010000",5,'1'); -- (2, 1, 2, 1, 2, 0, 0, 1, 0)
sync_reset;
check_mem(4247,"010100011","101010000",6,'1'); -- (2, 1, 2, 1, 2, 0, 0, 1, 1)
sync_reset;
check_mem(4248,"010100100","101010000",8,'1'); -- (2, 1, 2, 1, 2, 0, 1, 0, 0)
sync_reset;
check_mem(4249,"010100101","101010000",7,'1'); -- (2, 1, 2, 1, 2, 0, 1, 0, 1)
sync_reset;
check_mem(4250,"010100110","101010000",8,'1'); -- (2, 1, 2, 1, 2, 0, 1, 1, 0)
sync_reset;
check_mem(4251,"010100101","101010010",5,'1'); -- (2, 1, 2, 1, 2, 0, 1, 2, 1)
sync_reset;
check_mem(4252,"010101000","101010000",6,'1'); -- (2, 1, 2, 1, 2, 1, 0, 0, 0)
sync_reset;
check_mem(4253,"010101001","101010000",6,'1'); -- (2, 1, 2, 1, 2, 1, 0, 0, 1)
sync_reset;
check_mem(4254,"010101010","101010000",6,'1'); -- (2, 1, 2, 1, 2, 1, 0, 1, 0)
sync_reset;
check_mem(4255,"010101001","101010010",6,'1'); -- (2, 1, 2, 1, 2, 1, 0, 2, 1)
sync_reset;
check_mem(4256,"010101100","101010000",8,'1'); -- (2, 1, 2, 1, 2, 1, 1, 0, 0)
sync_reset;
check_mem(4257,"010101100","101010010",8,'1'); -- (2, 1, 2, 1, 2, 1, 1, 2, 0)
sync_reset;
check_mem(4258,"010100011","101011000",6,'1'); -- (2, 1, 2, 1, 2, 2, 0, 1, 1)
sync_reset;
check_mem(4259,"010100101","101011000",7,'1'); -- (2, 1, 2, 1, 2, 2, 1, 0, 1)
sync_reset;
check_mem(4260,"010100110","101011000",8,'1'); -- (2, 1, 2, 1, 2, 2, 1, 1, 0)
sync_reset;
check_mem(4261,"010000011","101100000",4,'1'); -- (2, 1, 2, 2, 0, 0, 0, 1, 1)
sync_reset;
check_mem(4262,"010000101","101100000",7,'1'); -- (2, 1, 2, 2, 0, 0, 1, 0, 1)
sync_reset;
check_mem(4263,"010000110","101100000",4,'1'); -- (2, 1, 2, 2, 0, 0, 1, 1, 0)
sync_reset;
check_mem(4264,"010001001","101100000",6,'1'); -- (2, 1, 2, 2, 0, 1, 0, 0, 1)
sync_reset;
check_mem(4265,"010001010","101100000",4,'1'); -- (2, 1, 2, 2, 0, 1, 0, 1, 0)
sync_reset;
check_mem(4266,"010001011","101100000",6,'1'); -- (2, 1, 2, 2, 0, 1, 0, 1, 1)
sync_reset;
check_mem(4267,"010001100","101100000",7,'1'); -- (2, 1, 2, 2, 0, 1, 1, 0, 0)
sync_reset;
check_mem(4268,"010001101","101100000",7,'1'); -- (2, 1, 2, 2, 0, 1, 1, 0, 1)
sync_reset;
check_mem(4269,"010001110","101100000",4,'1'); -- (2, 1, 2, 2, 0, 1, 1, 1, 0)
sync_reset;
check_mem(4270,"010001110","101100001",4,'1'); -- (2, 1, 2, 2, 0, 1, 1, 1, 2)
sync_reset;
check_mem(4271,"010001101","101100010",4,'1'); -- (2, 1, 2, 2, 0, 1, 1, 2, 1)
sync_reset;
check_mem(4272,"010010001","101100000",7,'1'); -- (2, 1, 2, 2, 1, 0, 0, 0, 1)
sync_reset;
check_mem(4273,"010010100","101100000",7,'1'); -- (2, 1, 2, 2, 1, 0, 1, 0, 0)
sync_reset;
check_mem(4274,"010010101","101100000",7,'1'); -- (2, 1, 2, 2, 1, 0, 1, 0, 1)
sync_reset;
check_mem(4275,"010010101","101100010",5,'1'); -- (2, 1, 2, 2, 1, 0, 1, 2, 1)
sync_reset;
check_mem(4276,"010011000","101100000",7,'1'); -- (2, 1, 2, 2, 1, 1, 0, 0, 0)
sync_reset;
check_mem(4277,"010011001","101100000",6,'1'); -- (2, 1, 2, 2, 1, 1, 0, 0, 1)
sync_reset;
check_mem(4278,"010011001","101100010",6,'1'); -- (2, 1, 2, 2, 1, 1, 0, 2, 1)
sync_reset;
check_mem(4279,"010011100","101100000",7,'1'); -- (2, 1, 2, 2, 1, 1, 1, 0, 0)
sync_reset;
check_mem(4280,"010011100","101100001",7,'1'); -- (2, 1, 2, 2, 1, 1, 1, 0, 2)
sync_reset;
check_mem(4281,"010011100","101100010",8,'1'); -- (2, 1, 2, 2, 1, 1, 1, 2, 0)
sync_reset;
check_mem(4282,"010010101","101101000",7,'1'); -- (2, 1, 2, 2, 1, 2, 1, 0, 1)
sync_reset;
check_mem(4283,"010001011","101110000",6,'1'); -- (2, 1, 2, 2, 2, 1, 0, 1, 1)
sync_reset;
check_mem(4284,"010001101","101110000",7,'1'); -- (2, 1, 2, 2, 2, 1, 1, 0, 1)
sync_reset;
check_mem(4285,"010001110","101110000",8,'1'); -- (2, 1, 2, 2, 2, 1, 1, 1, 0)
sync_reset;
check_mem(4286,"000000011","110000000",2,'1'); -- (2, 2, 0, 0, 0, 0, 0, 1, 1)
sync_reset;
check_mem(4287,"000000101","110000000",2,'1'); -- (2, 2, 0, 0, 0, 0, 1, 0, 1)
sync_reset;
check_mem(4288,"000000110","110000000",2,'1'); -- (2, 2, 0, 0, 0, 0, 1, 1, 0)
sync_reset;
check_mem(4289,"000001001","110000000",2,'1'); -- (2, 2, 0, 0, 0, 1, 0, 0, 1)
sync_reset;
check_mem(4290,"000001010","110000000",2,'1'); -- (2, 2, 0, 0, 0, 1, 0, 1, 0)
sync_reset;
check_mem(4291,"000001011","110000000",2,'1'); -- (2, 2, 0, 0, 0, 1, 0, 1, 1)
sync_reset;
check_mem(4292,"000001100","110000000",2,'1'); -- (2, 2, 0, 0, 0, 1, 1, 0, 0)
sync_reset;
check_mem(4293,"000001101","110000000",2,'1'); -- (2, 2, 0, 0, 0, 1, 1, 0, 1)
sync_reset;
check_mem(4294,"000001110","110000000",2,'1'); -- (2, 2, 0, 0, 0, 1, 1, 1, 0)
sync_reset;
check_mem(4295,"000001110","110000001",2,'1'); -- (2, 2, 0, 0, 0, 1, 1, 1, 2)
sync_reset;
check_mem(4296,"000001101","110000010",2,'1'); -- (2, 2, 0, 0, 0, 1, 1, 2, 1)
sync_reset;
check_mem(4297,"000001011","110000100",2,'1'); -- (2, 2, 0, 0, 0, 1, 2, 1, 1)
sync_reset;
check_mem(4298,"000010001","110000000",2,'1'); -- (2, 2, 0, 0, 1, 0, 0, 0, 1)
sync_reset;
check_mem(4299,"000010010","110000000",2,'1'); -- (2, 2, 0, 0, 1, 0, 0, 1, 0)
sync_reset;
check_mem(4300,"000010011","110000000",2,'1'); -- (2, 2, 0, 0, 1, 0, 0, 1, 1)
sync_reset;
check_mem(4301,"000010100","110000000",2,'1'); -- (2, 2, 0, 0, 1, 0, 1, 0, 0)
sync_reset;
check_mem(4302,"000010101","110000000",2,'1'); -- (2, 2, 0, 0, 1, 0, 1, 0, 1)
sync_reset;
check_mem(4303,"000010110","110000000",2,'1'); -- (2, 2, 0, 0, 1, 0, 1, 1, 0)
sync_reset;
check_mem(4304,"000010110","110000001",2,'1'); -- (2, 2, 0, 0, 1, 0, 1, 1, 2)
sync_reset;
check_mem(4305,"000010101","110000010",2,'1'); -- (2, 2, 0, 0, 1, 0, 1, 2, 1)
sync_reset;
check_mem(4306,"000010011","110000100",2,'1'); -- (2, 2, 0, 0, 1, 0, 2, 1, 1)
sync_reset;
check_mem(4307,"000011000","110000000",2,'1'); -- (2, 2, 0, 0, 1, 1, 0, 0, 0)
sync_reset;
check_mem(4308,"000011001","110000000",2,'1'); -- (2, 2, 0, 0, 1, 1, 0, 0, 1)
sync_reset;
check_mem(4309,"000011010","110000000",2,'1'); -- (2, 2, 0, 0, 1, 1, 0, 1, 0)
sync_reset;
check_mem(4310,"000011010","110000001",2,'1'); -- (2, 2, 0, 0, 1, 1, 0, 1, 2)
sync_reset;
check_mem(4311,"000011001","110000010",2,'1'); -- (2, 2, 0, 0, 1, 1, 0, 2, 1)
sync_reset;
check_mem(4312,"000011100","110000000",2,'1'); -- (2, 2, 0, 0, 1, 1, 1, 0, 0)
sync_reset;
check_mem(4313,"000011100","110000001",2,'1'); -- (2, 2, 0, 0, 1, 1, 1, 0, 2)
sync_reset;
check_mem(4314,"000011110","110000001",2,'1'); -- (2, 2, 0, 0, 1, 1, 1, 1, 2)
sync_reset;
check_mem(4315,"000011100","110000010",2,'1'); -- (2, 2, 0, 0, 1, 1, 1, 2, 0)
sync_reset;
check_mem(4316,"000011101","110000010",2,'1'); -- (2, 2, 0, 0, 1, 1, 1, 2, 1)
sync_reset;
check_mem(4317,"000011001","110000100",2,'1'); -- (2, 2, 0, 0, 1, 1, 2, 0, 1)
sync_reset;
check_mem(4318,"000011010","110000100",3,'1'); -- (2, 2, 0, 0, 1, 1, 2, 1, 0)
sync_reset;
check_mem(4319,"000011011","110000100",2,'1'); -- (2, 2, 0, 0, 1, 1, 2, 1, 1)
sync_reset;
check_mem(4320,"000010011","110001000",6,'1'); -- (2, 2, 0, 0, 1, 2, 0, 1, 1)
sync_reset;
check_mem(4321,"000010101","110001000",2,'1'); -- (2, 2, 0, 0, 1, 2, 1, 0, 1)
sync_reset;
check_mem(4322,"000010110","110001000",2,'1'); -- (2, 2, 0, 0, 1, 2, 1, 1, 0)
sync_reset;
check_mem(4323,"000001011","110010000",2,'1'); -- (2, 2, 0, 0, 2, 1, 0, 1, 1)
sync_reset;
check_mem(4324,"000001101","110010000",2,'1'); -- (2, 2, 0, 0, 2, 1, 1, 0, 1)
sync_reset;
check_mem(4325,"000001110","110010000",8,'1'); -- (2, 2, 0, 0, 2, 1, 1, 1, 0)
sync_reset;
check_mem(4326,"000100001","110000000",2,'1'); -- (2, 2, 0, 1, 0, 0, 0, 0, 1)
sync_reset;
check_mem(4327,"000100010","110000000",2,'1'); -- (2, 2, 0, 1, 0, 0, 0, 1, 0)
sync_reset;
check_mem(4328,"000100011","110000000",2,'1'); -- (2, 2, 0, 1, 0, 0, 0, 1, 1)
sync_reset;
check_mem(4329,"000100100","110000000",2,'1'); -- (2, 2, 0, 1, 0, 0, 1, 0, 0)
sync_reset;
check_mem(4330,"000100101","110000000",2,'1'); -- (2, 2, 0, 1, 0, 0, 1, 0, 1)
sync_reset;
check_mem(4331,"000100110","110000000",2,'1'); -- (2, 2, 0, 1, 0, 0, 1, 1, 0)
sync_reset;
check_mem(4332,"000100110","110000001",2,'1'); -- (2, 2, 0, 1, 0, 0, 1, 1, 2)
sync_reset;
check_mem(4333,"000100101","110000010",2,'1'); -- (2, 2, 0, 1, 0, 0, 1, 2, 1)
sync_reset;
check_mem(4334,"000100011","110000100",2,'1'); -- (2, 2, 0, 1, 0, 0, 2, 1, 1)
sync_reset;
check_mem(4335,"000101000","110000000",2,'1'); -- (2, 2, 0, 1, 0, 1, 0, 0, 0)
sync_reset;
check_mem(4336,"000101001","110000000",2,'1'); -- (2, 2, 0, 1, 0, 1, 0, 0, 1)
sync_reset;
check_mem(4337,"000101010","110000000",2,'1'); -- (2, 2, 0, 1, 0, 1, 0, 1, 0)
sync_reset;
check_mem(4338,"000101010","110000001",4,'1'); -- (2, 2, 0, 1, 0, 1, 0, 1, 2)
sync_reset;
check_mem(4339,"000101001","110000010",2,'1'); -- (2, 2, 0, 1, 0, 1, 0, 2, 1)
sync_reset;
check_mem(4340,"000101100","110000000",2,'1'); -- (2, 2, 0, 1, 0, 1, 1, 0, 0)
sync_reset;
check_mem(4341,"000101100","110000001",4,'1'); -- (2, 2, 0, 1, 0, 1, 1, 0, 2)
sync_reset;
check_mem(4342,"000101110","110000001",2,'1'); -- (2, 2, 0, 1, 0, 1, 1, 1, 2)
sync_reset;
check_mem(4343,"000101100","110000010",4,'1'); -- (2, 2, 0, 1, 0, 1, 1, 2, 0)
sync_reset;
check_mem(4344,"000101101","110000010",2,'1'); -- (2, 2, 0, 1, 0, 1, 1, 2, 1)
sync_reset;
check_mem(4345,"000101001","110000100",2,'1'); -- (2, 2, 0, 1, 0, 1, 2, 0, 1)
sync_reset;
check_mem(4346,"000101010","110000100",2,'1'); -- (2, 2, 0, 1, 0, 1, 2, 1, 0)
sync_reset;
check_mem(4347,"000101011","110000100",2,'1'); -- (2, 2, 0, 1, 0, 1, 2, 1, 1)
sync_reset;
check_mem(4348,"000100011","110001000",6,'1'); -- (2, 2, 0, 1, 0, 2, 0, 1, 1)
sync_reset;
check_mem(4349,"000100101","110001000",2,'1'); -- (2, 2, 0, 1, 0, 2, 1, 0, 1)
sync_reset;
check_mem(4350,"000100110","110001000",2,'1'); -- (2, 2, 0, 1, 0, 2, 1, 1, 0)
sync_reset;
check_mem(4351,"000110000","110000000",2,'1'); -- (2, 2, 0, 1, 1, 0, 0, 0, 0)
sync_reset;
check_mem(4352,"000110001","110000000",2,'1'); -- (2, 2, 0, 1, 1, 0, 0, 0, 1)
sync_reset;
check_mem(4353,"000110010","110000000",2,'1'); -- (2, 2, 0, 1, 1, 0, 0, 1, 0)
sync_reset;
check_mem(4354,"000110010","110000001",2,'1'); -- (2, 2, 0, 1, 1, 0, 0, 1, 2)
sync_reset;
check_mem(4355,"000110001","110000010",2,'1'); -- (2, 2, 0, 1, 1, 0, 0, 2, 1)
sync_reset;
check_mem(4356,"000110100","110000000",2,'1'); -- (2, 2, 0, 1, 1, 0, 1, 0, 0)
sync_reset;
check_mem(4357,"000110100","110000001",2,'1'); -- (2, 2, 0, 1, 1, 0, 1, 0, 2)
sync_reset;
check_mem(4358,"000110110","110000001",2,'1'); -- (2, 2, 0, 1, 1, 0, 1, 1, 2)
sync_reset;
check_mem(4359,"000110100","110000010",2,'1'); -- (2, 2, 0, 1, 1, 0, 1, 2, 0)
sync_reset;
check_mem(4360,"000110101","110000010",2,'1'); -- (2, 2, 0, 1, 1, 0, 1, 2, 1)
sync_reset;
check_mem(4361,"000110001","110000100",5,'1'); -- (2, 2, 0, 1, 1, 0, 2, 0, 1)
sync_reset;
check_mem(4362,"000110010","110000100",5,'1'); -- (2, 2, 0, 1, 1, 0, 2, 1, 0)
sync_reset;
check_mem(4363,"000110011","110000100",2,'1'); -- (2, 2, 0, 1, 1, 0, 2, 1, 1)
sync_reset;
check_mem(4364,"000110001","110001000",2,'1'); -- (2, 2, 0, 1, 1, 2, 0, 0, 1)
sync_reset;
check_mem(4365,"000110010","110001000",2,'1'); -- (2, 2, 0, 1, 1, 2, 0, 1, 0)
sync_reset;
check_mem(4366,"000110011","110001000",2,'1'); -- (2, 2, 0, 1, 1, 2, 0, 1, 1)
sync_reset;
check_mem(4367,"000110100","110001000",2,'1'); -- (2, 2, 0, 1, 1, 2, 1, 0, 0)
sync_reset;
check_mem(4368,"000110101","110001000",2,'1'); -- (2, 2, 0, 1, 1, 2, 1, 0, 1)
sync_reset;
check_mem(4369,"000110110","110001000",2,'1'); -- (2, 2, 0, 1, 1, 2, 1, 1, 0)
sync_reset;
check_mem(4370,"000110110","110001001",2,'1'); -- (2, 2, 0, 1, 1, 2, 1, 1, 2)
sync_reset;
check_mem(4371,"000110101","110001010",2,'1'); -- (2, 2, 0, 1, 1, 2, 1, 2, 1)
sync_reset;
check_mem(4372,"000110011","110001100",2,'1'); -- (2, 2, 0, 1, 1, 2, 2, 1, 1)
sync_reset;
check_mem(4373,"000100011","110010000",2,'1'); -- (2, 2, 0, 1, 2, 0, 0, 1, 1)
sync_reset;
check_mem(4374,"000100101","110010000",7,'1'); -- (2, 2, 0, 1, 2, 0, 1, 0, 1)
sync_reset;
check_mem(4375,"000100110","110010000",8,'1'); -- (2, 2, 0, 1, 2, 0, 1, 1, 0)
sync_reset;
check_mem(4376,"000101001","110010000",2,'1'); -- (2, 2, 0, 1, 2, 1, 0, 0, 1)
sync_reset;
check_mem(4377,"000101010","110010000",2,'1'); -- (2, 2, 0, 1, 2, 1, 0, 1, 0)
sync_reset;
check_mem(4378,"000101011","110010000",2,'1'); -- (2, 2, 0, 1, 2, 1, 0, 1, 1)
sync_reset;
check_mem(4379,"000101100","110010000",2,'1'); -- (2, 2, 0, 1, 2, 1, 1, 0, 0)
sync_reset;
check_mem(4380,"000101101","110010000",2,'1'); -- (2, 2, 0, 1, 2, 1, 1, 0, 1)
sync_reset;
check_mem(4381,"000101110","110010000",2,'1'); -- (2, 2, 0, 1, 2, 1, 1, 1, 0)
sync_reset;
check_mem(4382,"000101011","110010100",2,'1'); -- (2, 2, 0, 1, 2, 1, 2, 1, 1)
sync_reset;
check_mem(4383,"000001011","110100000",2,'1'); -- (2, 2, 0, 2, 0, 1, 0, 1, 1)
sync_reset;
check_mem(4384,"000001101","110100000",2,'1'); -- (2, 2, 0, 2, 0, 1, 1, 0, 1)
sync_reset;
check_mem(4385,"000001110","110100000",2,'1'); -- (2, 2, 0, 2, 0, 1, 1, 1, 0)
sync_reset;
check_mem(4386,"000010011","110100000",6,'1'); -- (2, 2, 0, 2, 1, 0, 0, 1, 1)
sync_reset;
check_mem(4387,"000010101","110100000",2,'1'); -- (2, 2, 0, 2, 1, 0, 1, 0, 1)
sync_reset;
check_mem(4388,"000010110","110100000",2,'1'); -- (2, 2, 0, 2, 1, 0, 1, 1, 0)
sync_reset;
check_mem(4389,"000011001","110100000",2,'1'); -- (2, 2, 0, 2, 1, 1, 0, 0, 1)
sync_reset;
check_mem(4390,"000011010","110100000",2,'1'); -- (2, 2, 0, 2, 1, 1, 0, 1, 0)
sync_reset;
check_mem(4391,"000011011","110100000",2,'1'); -- (2, 2, 0, 2, 1, 1, 0, 1, 1)
sync_reset;
check_mem(4392,"000011100","110100000",2,'1'); -- (2, 2, 0, 2, 1, 1, 1, 0, 0)
sync_reset;
check_mem(4393,"000011101","110100000",2,'1'); -- (2, 2, 0, 2, 1, 1, 1, 0, 1)
sync_reset;
check_mem(4394,"000011110","110100000",2,'1'); -- (2, 2, 0, 2, 1, 1, 1, 1, 0)
sync_reset;
check_mem(4395,"000011110","110100001",2,'1'); -- (2, 2, 0, 2, 1, 1, 1, 1, 2)
sync_reset;
check_mem(4396,"000011101","110100010",2,'1'); -- (2, 2, 0, 2, 1, 1, 1, 2, 1)
sync_reset;
check_mem(4397,"001000001","110000000",3,'1'); -- (2, 2, 1, 0, 0, 0, 0, 0, 1)
sync_reset;
check_mem(4398,"001000010","110000000",3,'1'); -- (2, 2, 1, 0, 0, 0, 0, 1, 0)
sync_reset;
check_mem(4399,"001000011","110000000",3,'1'); -- (2, 2, 1, 0, 0, 0, 0, 1, 1)
sync_reset;
check_mem(4400,"001000100","110000000",4,'1'); -- (2, 2, 1, 0, 0, 0, 1, 0, 0)
sync_reset;
check_mem(4401,"001000101","110000000",3,'1'); -- (2, 2, 1, 0, 0, 0, 1, 0, 1)
sync_reset;
check_mem(4402,"001000110","110000000",3,'1'); -- (2, 2, 1, 0, 0, 0, 1, 1, 0)
sync_reset;
check_mem(4403,"001000110","110000001",4,'1'); -- (2, 2, 1, 0, 0, 0, 1, 1, 2)
sync_reset;
check_mem(4404,"001000101","110000010",4,'1'); -- (2, 2, 1, 0, 0, 0, 1, 2, 1)
sync_reset;
check_mem(4405,"001000011","110000100",5,'1'); -- (2, 2, 1, 0, 0, 0, 2, 1, 1)
sync_reset;
check_mem(4406,"001001000","110000000",3,'1'); -- (2, 2, 1, 0, 0, 1, 0, 0, 0)
sync_reset;
check_mem(4407,"001001010","110000000",3,'1'); -- (2, 2, 1, 0, 0, 1, 0, 1, 0)
sync_reset;
check_mem(4408,"001001010","110000001",4,'1'); -- (2, 2, 1, 0, 0, 1, 0, 1, 2)
sync_reset;
check_mem(4409,"001001100","110000000",3,'1'); -- (2, 2, 1, 0, 0, 1, 1, 0, 0)
sync_reset;
check_mem(4410,"001001100","110000001",4,'1'); -- (2, 2, 1, 0, 0, 1, 1, 0, 2)
sync_reset;
check_mem(4411,"001001110","110000001",4,'1'); -- (2, 2, 1, 0, 0, 1, 1, 1, 2)
sync_reset;
check_mem(4412,"001001100","110000010",4,'1'); -- (2, 2, 1, 0, 0, 1, 1, 2, 0)
sync_reset;
check_mem(4413,"001001010","110000100",3,'1'); -- (2, 2, 1, 0, 0, 1, 2, 1, 0)
sync_reset;
check_mem(4414,"001000011","110001000",6,'1'); -- (2, 2, 1, 0, 0, 2, 0, 1, 1)
sync_reset;
check_mem(4415,"001000101","110001000",3,'1'); -- (2, 2, 1, 0, 0, 2, 1, 0, 1)
sync_reset;
check_mem(4416,"001000110","110001000",3,'1'); -- (2, 2, 1, 0, 0, 2, 1, 1, 0)
sync_reset;
check_mem(4417,"001010000","110000000",3,'1'); -- (2, 2, 1, 0, 1, 0, 0, 0, 0)
sync_reset;
check_mem(4418,"001010001","110000000",3,'1'); -- (2, 2, 1, 0, 1, 0, 0, 0, 1)
sync_reset;
check_mem(4419,"001010010","110000000",6,'1'); -- (2, 2, 1, 0, 1, 0, 0, 1, 0)
sync_reset;
check_mem(4420,"001010010","110000001",3,'1'); -- (2, 2, 1, 0, 1, 0, 0, 1, 2)
sync_reset;
check_mem(4421,"001010001","110000010",3,'1'); -- (2, 2, 1, 0, 1, 0, 0, 2, 1)
sync_reset;
check_mem(4422,"001010001","110000100",5,'1'); -- (2, 2, 1, 0, 1, 0, 2, 0, 1)
sync_reset;
check_mem(4423,"001010010","110000100",3,'1'); -- (2, 2, 1, 0, 1, 0, 2, 1, 0)
sync_reset;
check_mem(4424,"001010011","110000100",3,'1'); -- (2, 2, 1, 0, 1, 0, 2, 1, 1)
sync_reset;
check_mem(4425,"001011000","110000000",3,'1'); -- (2, 2, 1, 0, 1, 1, 0, 0, 0)
sync_reset;
check_mem(4426,"001011000","110000001",3,'1'); -- (2, 2, 1, 0, 1, 1, 0, 0, 2)
sync_reset;
check_mem(4427,"001011010","110000001",3,'1'); -- (2, 2, 1, 0, 1, 1, 0, 1, 2)
sync_reset;
check_mem(4428,"001011000","110000010",3,'1'); -- (2, 2, 1, 0, 1, 1, 0, 2, 0)
sync_reset;
check_mem(4429,"001011000","110000100",3,'1'); -- (2, 2, 1, 0, 1, 1, 2, 0, 0)
sync_reset;
check_mem(4430,"001011010","110000100",3,'1'); -- (2, 2, 1, 0, 1, 1, 2, 1, 0)
sync_reset;
check_mem(4431,"001011010","110000101",3,'1'); -- (2, 2, 1, 0, 1, 1, 2, 1, 2)
sync_reset;
check_mem(4432,"001010001","110001000",6,'1'); -- (2, 2, 1, 0, 1, 2, 0, 0, 1)
sync_reset;
check_mem(4433,"001010010","110001000",6,'1'); -- (2, 2, 1, 0, 1, 2, 0, 1, 0)
sync_reset;
check_mem(4434,"001010011","110001000",6,'1'); -- (2, 2, 1, 0, 1, 2, 0, 1, 1)
sync_reset;
check_mem(4435,"001010011","110001100",3,'1'); -- (2, 2, 1, 0, 1, 2, 2, 1, 1)
sync_reset;
check_mem(4436,"001000011","110010000",3,'1'); -- (2, 2, 1, 0, 2, 0, 0, 1, 1)
sync_reset;
check_mem(4437,"001000101","110010000",5,'1'); -- (2, 2, 1, 0, 2, 0, 1, 0, 1)
sync_reset;
check_mem(4438,"001000110","110010000",8,'1'); -- (2, 2, 1, 0, 2, 0, 1, 1, 0)
sync_reset;
check_mem(4439,"001001010","110010000",8,'1'); -- (2, 2, 1, 0, 2, 1, 0, 1, 0)
sync_reset;
check_mem(4440,"001001100","110010000",8,'1'); -- (2, 2, 1, 0, 2, 1, 1, 0, 0)
sync_reset;
check_mem(4441,"001001110","110010000",8,'1'); -- (2, 2, 1, 0, 2, 1, 1, 1, 0)
sync_reset;
check_mem(4442,"001100000","110000000",4,'1'); -- (2, 2, 1, 1, 0, 0, 0, 0, 0)
sync_reset;
check_mem(4443,"001100001","110000000",4,'1'); -- (2, 2, 1, 1, 0, 0, 0, 0, 1)
sync_reset;
check_mem(4444,"001100010","110000000",4,'1'); -- (2, 2, 1, 1, 0, 0, 0, 1, 0)
sync_reset;
check_mem(4445,"001100010","110000001",4,'1'); -- (2, 2, 1, 1, 0, 0, 0, 1, 2)
sync_reset;
check_mem(4446,"001100001","110000010",4,'1'); -- (2, 2, 1, 1, 0, 0, 0, 2, 1)
sync_reset;
check_mem(4447,"001100100","110000000",4,'1'); -- (2, 2, 1, 1, 0, 0, 1, 0, 0)
sync_reset;
check_mem(4448,"001100100","110000001",4,'1'); -- (2, 2, 1, 1, 0, 0, 1, 0, 2)
sync_reset;
check_mem(4449,"001100110","110000001",4,'1'); -- (2, 2, 1, 1, 0, 0, 1, 1, 2)
sync_reset;
check_mem(4450,"001100100","110000010",4,'1'); -- (2, 2, 1, 1, 0, 0, 1, 2, 0)
sync_reset;
check_mem(4451,"001100101","110000010",4,'1'); -- (2, 2, 1, 1, 0, 0, 1, 2, 1)
sync_reset;
check_mem(4452,"001100001","110000100",5,'1'); -- (2, 2, 1, 1, 0, 0, 2, 0, 1)
sync_reset;
check_mem(4453,"001100010","110000100",5,'1'); -- (2, 2, 1, 1, 0, 0, 2, 1, 0)
sync_reset;
check_mem(4454,"001100011","110000100",5,'1'); -- (2, 2, 1, 1, 0, 0, 2, 1, 1)
sync_reset;
check_mem(4455,"001101000","110000000",4,'1'); -- (2, 2, 1, 1, 0, 1, 0, 0, 0)
sync_reset;
check_mem(4456,"001101000","110000001",4,'1'); -- (2, 2, 1, 1, 0, 1, 0, 0, 2)
sync_reset;
check_mem(4457,"001101010","110000001",4,'1'); -- (2, 2, 1, 1, 0, 1, 0, 1, 2)
sync_reset;
check_mem(4458,"001101000","110000010",4,'1'); -- (2, 2, 1, 1, 0, 1, 0, 2, 0)
sync_reset;
check_mem(4459,"001101100","110000001",4,'1'); -- (2, 2, 1, 1, 0, 1, 1, 0, 2)
sync_reset;
check_mem(4460,"001101100","110000010",4,'1'); -- (2, 2, 1, 1, 0, 1, 1, 2, 0)
sync_reset;
check_mem(4461,"001101100","110000011",4,'1'); -- (2, 2, 1, 1, 0, 1, 1, 2, 2)
sync_reset;
check_mem(4462,"001101000","110000100",4,'1'); -- (2, 2, 1, 1, 0, 1, 2, 0, 0)
sync_reset;
check_mem(4463,"001101010","110000100",4,'1'); -- (2, 2, 1, 1, 0, 1, 2, 1, 0)
sync_reset;
check_mem(4464,"001101010","110000101",4,'1'); -- (2, 2, 1, 1, 0, 1, 2, 1, 2)
sync_reset;
check_mem(4465,"001100001","110001000",6,'1'); -- (2, 2, 1, 1, 0, 2, 0, 0, 1)
sync_reset;
check_mem(4466,"001100010","110001000",6,'1'); -- (2, 2, 1, 1, 0, 2, 0, 1, 0)
sync_reset;
check_mem(4467,"001100011","110001000",6,'1'); -- (2, 2, 1, 1, 0, 2, 0, 1, 1)
sync_reset;
check_mem(4468,"001100100","110001000",4,'1'); -- (2, 2, 1, 1, 0, 2, 1, 0, 0)
sync_reset;
check_mem(4469,"001100101","110001000",4,'1'); -- (2, 2, 1, 1, 0, 2, 1, 0, 1)
sync_reset;
check_mem(4470,"001100110","110001000",4,'1'); -- (2, 2, 1, 1, 0, 2, 1, 1, 0)
sync_reset;
check_mem(4471,"001100110","110001001",4,'1'); -- (2, 2, 1, 1, 0, 2, 1, 1, 2)
sync_reset;
check_mem(4472,"001100101","110001010",4,'1'); -- (2, 2, 1, 1, 0, 2, 1, 2, 1)
sync_reset;
check_mem(4473,"001100011","110001100",4,'1'); -- (2, 2, 1, 1, 0, 2, 2, 1, 1)
sync_reset;
check_mem(4474,"001110000","110000000",5,'1'); -- (2, 2, 1, 1, 1, 0, 0, 0, 0)
sync_reset;
check_mem(4475,"001110000","110000001",5,'1'); -- (2, 2, 1, 1, 1, 0, 0, 0, 2)
sync_reset;
check_mem(4476,"001110010","110000001",5,'1'); -- (2, 2, 1, 1, 1, 0, 0, 1, 2)
sync_reset;
check_mem(4477,"001110000","110000010",5,'1'); -- (2, 2, 1, 1, 1, 0, 0, 2, 0)
sync_reset;
check_mem(4478,"001110001","110000010",5,'1'); -- (2, 2, 1, 1, 1, 0, 0, 2, 1)
sync_reset;
check_mem(4479,"001110000","110000100",5,'1'); -- (2, 2, 1, 1, 1, 0, 2, 0, 0)
sync_reset;
check_mem(4480,"001110001","110000100",5,'1'); -- (2, 2, 1, 1, 1, 0, 2, 0, 1)
sync_reset;
check_mem(4481,"001110010","110000100",5,'1'); -- (2, 2, 1, 1, 1, 0, 2, 1, 0)
sync_reset;
check_mem(4482,"001110010","110000101",5,'1'); -- (2, 2, 1, 1, 1, 0, 2, 1, 2)
sync_reset;
check_mem(4483,"001110001","110000110",5,'1'); -- (2, 2, 1, 1, 1, 0, 2, 2, 1)
sync_reset;
check_mem(4484,"001110000","110001000",6,'1'); -- (2, 2, 1, 1, 1, 2, 0, 0, 0)
sync_reset;
check_mem(4485,"001110001","110001000",6,'1'); -- (2, 2, 1, 1, 1, 2, 0, 0, 1)
sync_reset;
check_mem(4486,"001110010","110001000",6,'1'); -- (2, 2, 1, 1, 1, 2, 0, 1, 0)
sync_reset;
check_mem(4487,"001110010","110001001",6,'1'); -- (2, 2, 1, 1, 1, 2, 0, 1, 2)
sync_reset;
check_mem(4488,"001110001","110001010",6,'1'); -- (2, 2, 1, 1, 1, 2, 0, 2, 1)
sync_reset;
check_mem(4489,"001110001","110001100",7,'1'); -- (2, 2, 1, 1, 1, 2, 2, 0, 1)
sync_reset;
check_mem(4490,"001110010","110001100",8,'1'); -- (2, 2, 1, 1, 1, 2, 2, 1, 0)
sync_reset;
check_mem(4491,"001100001","110010000",5,'1'); -- (2, 2, 1, 1, 2, 0, 0, 0, 1)
sync_reset;
check_mem(4492,"001100010","110010000",8,'1'); -- (2, 2, 1, 1, 2, 0, 0, 1, 0)
sync_reset;
check_mem(4493,"001100011","110010000",5,'1'); -- (2, 2, 1, 1, 2, 0, 0, 1, 1)
sync_reset;
check_mem(4494,"001100100","110010000",5,'1'); -- (2, 2, 1, 1, 2, 0, 1, 0, 0)
sync_reset;
check_mem(4495,"001100101","110010000",7,'1'); -- (2, 2, 1, 1, 2, 0, 1, 0, 1)
sync_reset;
check_mem(4496,"001100110","110010000",8,'1'); -- (2, 2, 1, 1, 2, 0, 1, 1, 0)
sync_reset;
check_mem(4497,"001100011","110010100",5,'1'); -- (2, 2, 1, 1, 2, 0, 2, 1, 1)
sync_reset;
check_mem(4498,"001101000","110010000",8,'1'); -- (2, 2, 1, 1, 2, 1, 0, 0, 0)
sync_reset;
check_mem(4499,"001101010","110010000",8,'1'); -- (2, 2, 1, 1, 2, 1, 0, 1, 0)
sync_reset;
check_mem(4500,"001101100","110010000",7,'1'); -- (2, 2, 1, 1, 2, 1, 1, 0, 0)
sync_reset;
check_mem(4501,"001101010","110010100",8,'1'); -- (2, 2, 1, 1, 2, 1, 2, 1, 0)
sync_reset;
check_mem(4502,"001100011","110011000",6,'1'); -- (2, 2, 1, 1, 2, 2, 0, 1, 1)
sync_reset;
check_mem(4503,"001100101","110011000",7,'1'); -- (2, 2, 1, 1, 2, 2, 1, 0, 1)
sync_reset;
check_mem(4504,"001100110","110011000",8,'1'); -- (2, 2, 1, 1, 2, 2, 1, 1, 0)
sync_reset;
check_mem(4505,"001000011","110100000",5,'1'); -- (2, 2, 1, 2, 0, 0, 0, 1, 1)
sync_reset;
check_mem(4506,"001000101","110100000",4,'1'); -- (2, 2, 1, 2, 0, 0, 1, 0, 1)
sync_reset;
check_mem(4507,"001000110","110100000",4,'1'); -- (2, 2, 1, 2, 0, 0, 1, 1, 0)
sync_reset;
check_mem(4508,"001001010","110100000",6,'1'); -- (2, 2, 1, 2, 0, 1, 0, 1, 0)
sync_reset;
check_mem(4509,"001001100","110100000",4,'1'); -- (2, 2, 1, 2, 0, 1, 1, 0, 0)
sync_reset;
check_mem(4510,"001001110","110100000",4,'1'); -- (2, 2, 1, 2, 0, 1, 1, 1, 0)
sync_reset;
check_mem(4511,"001001110","110100001",4,'1'); -- (2, 2, 1, 2, 0, 1, 1, 1, 2)
sync_reset;
check_mem(4512,"001010001","110100000",5,'1'); -- (2, 2, 1, 2, 1, 0, 0, 0, 1)
sync_reset;
check_mem(4513,"001010010","110100000",6,'1'); -- (2, 2, 1, 2, 1, 0, 0, 1, 0)
sync_reset;
check_mem(4514,"001010011","110100000",6,'1'); -- (2, 2, 1, 2, 1, 0, 0, 1, 1)
sync_reset;
check_mem(4515,"001011000","110100000",6,'1'); -- (2, 2, 1, 2, 1, 1, 0, 0, 0)
sync_reset;
check_mem(4516,"001011010","110100000",6,'1'); -- (2, 2, 1, 2, 1, 1, 0, 1, 0)
sync_reset;
check_mem(4517,"001011010","110100001",6,'1'); -- (2, 2, 1, 2, 1, 1, 0, 1, 2)
sync_reset;
check_mem(4518,"001010011","110101000",6,'1'); -- (2, 2, 1, 2, 1, 2, 0, 1, 1)
sync_reset;
check_mem(4519,"001001110","110110000",8,'1'); -- (2, 2, 1, 2, 2, 1, 1, 1, 0)
--
-- Some non-matching cases

sync_reset;
check_mem(4519,"001111110","110111100",8,'0');
sync_reset;
check_mem(2874,"100111011","010001101",4,'0'); -- (1, 2, 0, 1, 0, 2, 2, 1, 1)
sync_reset;
check_mem(251,"000001010","000110001",8,'0'); -- (0, 0, 0, 2, 2, 1, 0, 1, 0)
sync_reset;
check_mem(4518,"001011010","110100001",6,'0'); -- (2, 2, 1, 2, 1, 1, 0, 1, 2)

		report "#### TESTS COMPLETED ####";
        sim_finished <= true;
        wait;
        
    end process simulation;


end test;
